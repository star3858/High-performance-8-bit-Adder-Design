magic
tech tsmc
timestamp 1513082383
<< nwell >>
rect -2783 925 117 957
rect -672 924 -656 925
rect -3105 593 -1750 625
rect -1674 591 -81 623
rect -71 591 96 623
rect -2847 369 87 402
<< ntransistor >>
rect -2765 811 -2762 819
rect -2694 822 -2691 830
rect -2678 822 -2675 830
rect -2662 822 -2659 830
rect -2645 822 -2642 830
rect -2723 810 -2720 818
rect -2609 796 -2606 804
rect -2593 796 -2590 804
rect -2565 796 -2562 804
rect -2312 811 -2309 819
rect -2241 822 -2238 830
rect -2225 822 -2222 830
rect -2209 822 -2206 830
rect -2192 822 -2189 830
rect -2270 810 -2267 818
rect -2156 796 -2153 804
rect -2140 796 -2137 804
rect -2112 796 -2109 804
rect -2021 811 -2018 819
rect -1950 822 -1947 830
rect -1934 822 -1931 830
rect -1918 822 -1915 830
rect -1901 822 -1898 830
rect -1979 810 -1976 818
rect -1865 796 -1862 804
rect -1849 796 -1846 804
rect -1821 796 -1818 804
rect -1778 811 -1775 819
rect -1707 822 -1704 830
rect -1691 822 -1688 830
rect -1675 822 -1672 830
rect -1658 822 -1655 830
rect -1736 810 -1733 818
rect -1622 796 -1619 804
rect -1606 796 -1603 804
rect -1578 796 -1575 804
rect -1096 811 -1093 819
rect -1025 822 -1022 830
rect -1009 822 -1006 830
rect -993 822 -990 830
rect -976 822 -973 830
rect -1054 810 -1051 818
rect -940 796 -937 804
rect -924 796 -921 804
rect -896 796 -893 804
rect -643 811 -640 819
rect -572 822 -569 830
rect -556 822 -553 830
rect -540 822 -537 830
rect -523 822 -520 830
rect -601 810 -598 818
rect -3087 483 -3084 491
rect -3070 483 -3067 491
rect -3054 483 -3051 491
rect -3038 483 -3035 491
rect -3022 483 -3019 491
rect -2994 483 -2991 491
rect -2959 483 -2956 491
rect -2943 483 -2940 491
rect -2927 483 -2924 491
rect -2911 483 -2908 491
rect -2883 483 -2880 491
rect -2850 483 -2847 491
rect -2834 483 -2831 491
rect -2818 483 -2815 491
rect -2790 483 -2787 491
rect -2751 483 -2748 491
rect -2735 483 -2732 491
rect -2707 483 -2704 491
rect -2673 483 -2670 491
rect -2657 483 -2654 491
rect -2641 483 -2638 491
rect -2625 483 -2622 491
rect -2610 483 -2607 491
rect -2582 483 -2579 491
rect -2516 483 -2513 491
rect -2500 483 -2497 491
rect -2484 483 -2481 491
rect -2468 483 -2465 491
rect -2440 483 -2437 491
rect -2407 483 -2404 491
rect -2391 483 -2388 491
rect -2375 483 -2372 491
rect -2347 483 -2344 491
rect -2308 483 -2305 491
rect -2292 483 -2289 491
rect -2264 483 -2261 491
rect -2230 483 -2227 491
rect -2214 483 -2211 491
rect -2198 483 -2195 491
rect -2182 483 -2179 491
rect -2154 483 -2151 491
rect -2033 483 -2030 491
rect -2017 483 -2014 491
rect -2001 483 -1998 491
rect -1973 483 -1970 491
rect -1934 483 -1931 491
rect -1918 483 -1915 491
rect -1890 483 -1887 491
rect -1833 483 -1830 491
rect -1817 483 -1814 491
rect -1800 483 -1797 491
rect -1772 483 -1769 491
rect -1653 481 -1650 489
rect -1637 481 -1634 489
rect -1609 481 -1606 489
rect -1574 481 -1571 489
rect -1557 481 -1554 489
rect -1529 481 -1526 489
rect -2829 274 -2826 282
rect -2761 285 -2758 293
rect -2745 285 -2742 293
rect -2729 285 -2726 293
rect -2713 285 -2710 293
rect -2790 273 -2787 281
rect -487 796 -484 804
rect -471 796 -468 804
rect -443 796 -440 804
rect -352 811 -349 819
rect -281 822 -278 830
rect -265 822 -262 830
rect -249 822 -246 830
rect -232 822 -229 830
rect -310 810 -307 818
rect -196 796 -193 804
rect -180 796 -177 804
rect -152 796 -149 804
rect -109 811 -106 819
rect -38 822 -35 830
rect -22 822 -19 830
rect -6 822 -3 830
rect 11 822 14 830
rect -67 810 -64 818
rect 47 796 50 804
rect 63 796 66 804
rect 91 796 94 804
rect -1483 481 -1480 489
rect -1466 481 -1463 489
rect -1450 481 -1447 489
rect -1434 481 -1431 489
rect -1418 481 -1415 489
rect -1390 481 -1387 489
rect -1355 481 -1352 489
rect -1339 481 -1336 489
rect -1323 481 -1320 489
rect -1307 481 -1304 489
rect -1279 481 -1276 489
rect -1246 481 -1243 489
rect -1230 481 -1227 489
rect -1214 481 -1211 489
rect -1186 481 -1183 489
rect -1147 481 -1144 489
rect -1131 481 -1128 489
rect -1103 481 -1100 489
rect -1069 481 -1066 489
rect -1053 481 -1050 489
rect -1037 481 -1034 489
rect -1021 481 -1018 489
rect -1006 481 -1003 489
rect -978 481 -975 489
rect -847 481 -844 489
rect -831 481 -828 489
rect -815 481 -812 489
rect -799 481 -796 489
rect -771 481 -768 489
rect -738 481 -735 489
rect -722 481 -719 489
rect -706 481 -703 489
rect -678 481 -675 489
rect -639 481 -636 489
rect -623 481 -620 489
rect -595 481 -592 489
rect -561 481 -558 489
rect -545 481 -542 489
rect -529 481 -526 489
rect -513 481 -510 489
rect -485 481 -482 489
rect -2321 274 -2318 282
rect -2253 285 -2250 293
rect -2237 285 -2234 293
rect -2221 285 -2218 293
rect -2205 285 -2202 293
rect -2282 273 -2279 281
rect -1977 274 -1974 282
rect -1909 285 -1906 293
rect -1893 285 -1890 293
rect -1877 285 -1874 293
rect -1861 285 -1858 293
rect -1938 273 -1935 281
rect -364 481 -361 489
rect -348 481 -345 489
rect -332 481 -329 489
rect -304 481 -301 489
rect -265 481 -262 489
rect -249 481 -246 489
rect -221 481 -218 489
rect -164 481 -161 489
rect -148 481 -145 489
rect -131 481 -128 489
rect -103 481 -100 489
rect -50 481 -47 489
rect -34 481 -31 489
rect -6 481 -3 489
rect 29 481 32 489
rect 46 481 49 489
rect 74 481 77 489
rect -1596 274 -1593 282
rect -1528 285 -1525 293
rect -1512 285 -1509 293
rect -1496 285 -1493 293
rect -1480 285 -1477 293
rect -1557 273 -1554 281
rect -1160 274 -1157 282
rect -1092 285 -1089 293
rect -1076 285 -1073 293
rect -1060 285 -1057 293
rect -1044 285 -1041 293
rect -1121 273 -1118 281
rect -652 274 -649 282
rect -584 285 -581 293
rect -568 285 -565 293
rect -552 285 -549 293
rect -536 285 -533 293
rect -613 273 -610 281
rect -308 274 -305 282
rect -240 285 -237 293
rect -224 285 -221 293
rect -208 285 -205 293
rect -192 285 -189 293
rect -269 273 -266 281
rect -50 274 -47 282
rect 18 285 21 293
rect 34 285 37 293
rect 50 285 53 293
rect 66 285 69 293
rect -11 273 -8 281
<< ptransistor >>
rect -2765 933 -2762 949
rect -2723 933 -2720 949
rect -2694 933 -2691 949
rect -2678 933 -2675 949
rect -2662 933 -2659 949
rect -2645 933 -2642 949
rect -2609 933 -2606 949
rect -2593 933 -2590 949
rect -2565 933 -2562 949
rect -2312 933 -2309 949
rect -2270 933 -2267 949
rect -2241 933 -2238 949
rect -2225 933 -2222 949
rect -2209 933 -2206 949
rect -2192 933 -2189 949
rect -2156 933 -2153 949
rect -2140 933 -2137 949
rect -2112 933 -2109 949
rect -2021 933 -2018 949
rect -1979 933 -1976 949
rect -1950 933 -1947 949
rect -1934 933 -1931 949
rect -1918 933 -1915 949
rect -1901 933 -1898 949
rect -1865 933 -1862 949
rect -1849 933 -1846 949
rect -1821 933 -1818 949
rect -1778 933 -1775 949
rect -1736 933 -1733 949
rect -1707 933 -1704 949
rect -1691 933 -1688 949
rect -1675 933 -1672 949
rect -1658 933 -1655 949
rect -1622 933 -1619 949
rect -1606 933 -1603 949
rect -1578 933 -1575 949
rect -1096 933 -1093 949
rect -1054 933 -1051 949
rect -1025 933 -1022 949
rect -1009 933 -1006 949
rect -993 933 -990 949
rect -976 933 -973 949
rect -940 933 -937 949
rect -924 933 -921 949
rect -896 933 -893 949
rect -643 933 -640 949
rect -601 933 -598 949
rect -572 933 -569 949
rect -556 933 -553 949
rect -540 933 -537 949
rect -523 933 -520 949
rect -487 933 -484 949
rect -471 933 -468 949
rect -443 933 -440 949
rect -352 933 -349 949
rect -310 933 -307 949
rect -281 933 -278 949
rect -265 933 -262 949
rect -249 933 -246 949
rect -232 933 -229 949
rect -196 933 -193 949
rect -180 933 -177 949
rect -152 933 -149 949
rect -109 933 -106 949
rect -67 933 -64 949
rect -38 933 -35 949
rect -22 933 -19 949
rect -6 933 -3 949
rect 11 933 14 949
rect 47 933 50 949
rect 63 933 66 949
rect 91 933 94 949
rect -3087 601 -3084 617
rect -3070 601 -3067 617
rect -3054 601 -3051 617
rect -3038 601 -3035 617
rect -3022 601 -3019 617
rect -2994 601 -2991 617
rect -2959 601 -2956 617
rect -2943 601 -2940 617
rect -2927 601 -2924 617
rect -2911 601 -2908 617
rect -2883 601 -2880 617
rect -2850 601 -2847 617
rect -2834 601 -2831 617
rect -2818 601 -2815 617
rect -2790 601 -2787 617
rect -2751 601 -2748 617
rect -2735 601 -2732 617
rect -2707 601 -2704 617
rect -2673 601 -2670 617
rect -2657 601 -2654 617
rect -2641 601 -2638 617
rect -2625 601 -2622 617
rect -2610 601 -2607 617
rect -2582 601 -2579 617
rect -2516 601 -2513 617
rect -2500 601 -2497 617
rect -2484 601 -2481 617
rect -2468 601 -2465 617
rect -2440 601 -2437 617
rect -2407 601 -2404 617
rect -2391 601 -2388 617
rect -2375 601 -2372 617
rect -2347 601 -2344 617
rect -2308 601 -2305 617
rect -2292 601 -2289 617
rect -2264 601 -2261 617
rect -2230 601 -2227 617
rect -2214 601 -2211 617
rect -2198 601 -2195 617
rect -2182 601 -2179 617
rect -2154 601 -2151 617
rect -2033 601 -2030 617
rect -2017 601 -2014 617
rect -2001 601 -1998 617
rect -1973 601 -1970 617
rect -1934 601 -1931 617
rect -1918 601 -1915 617
rect -1890 601 -1887 617
rect -1833 601 -1830 617
rect -1817 601 -1814 617
rect -1800 601 -1797 617
rect -1772 601 -1769 617
rect -2829 378 -2826 394
rect -2790 378 -2787 394
rect -1653 599 -1650 615
rect -1637 599 -1634 615
rect -1609 599 -1606 615
rect -1574 599 -1571 615
rect -1557 599 -1554 615
rect -1529 599 -1526 615
rect -1483 599 -1480 615
rect -1466 599 -1463 615
rect -1450 599 -1447 615
rect -1434 599 -1431 615
rect -1418 599 -1415 615
rect -1390 599 -1387 615
rect -1355 599 -1352 615
rect -1339 599 -1336 615
rect -1323 599 -1320 615
rect -1307 599 -1304 615
rect -1279 599 -1276 615
rect -1246 599 -1243 615
rect -1230 599 -1227 615
rect -1214 599 -1211 615
rect -1186 599 -1183 615
rect -1147 599 -1144 615
rect -1131 599 -1128 615
rect -1103 599 -1100 615
rect -1069 599 -1066 615
rect -1053 599 -1050 615
rect -1037 599 -1034 615
rect -1021 599 -1018 615
rect -1006 599 -1003 615
rect -978 599 -975 615
rect -2761 377 -2758 393
rect -2745 377 -2742 393
rect -2729 377 -2726 393
rect -2713 377 -2710 393
rect -2321 378 -2318 394
rect -2282 378 -2279 394
rect -2253 377 -2250 393
rect -2237 377 -2234 393
rect -2221 377 -2218 393
rect -2205 377 -2202 393
rect -1977 378 -1974 394
rect -1938 378 -1935 394
rect -847 599 -844 615
rect -831 599 -828 615
rect -815 599 -812 615
rect -799 599 -796 615
rect -771 599 -768 615
rect -738 599 -735 615
rect -722 599 -719 615
rect -706 599 -703 615
rect -678 599 -675 615
rect -639 599 -636 615
rect -623 599 -620 615
rect -595 599 -592 615
rect -561 599 -558 615
rect -545 599 -542 615
rect -529 599 -526 615
rect -513 599 -510 615
rect -485 599 -482 615
rect -364 599 -361 615
rect -348 599 -345 615
rect -332 599 -329 615
rect -304 599 -301 615
rect -265 599 -262 615
rect -249 599 -246 615
rect -221 599 -218 615
rect -164 599 -161 615
rect -148 599 -145 615
rect -131 599 -128 615
rect -103 599 -100 615
rect -50 599 -47 615
rect -34 599 -31 615
rect -6 599 -3 615
rect 29 599 32 615
rect 46 599 49 615
rect 74 599 77 615
rect -1909 377 -1906 393
rect -1893 377 -1890 393
rect -1877 377 -1874 393
rect -1861 377 -1858 393
rect -1596 378 -1593 394
rect -1557 378 -1554 394
rect -1528 377 -1525 393
rect -1512 377 -1509 393
rect -1496 377 -1493 393
rect -1480 377 -1477 393
rect -1160 378 -1157 394
rect -1121 378 -1118 394
rect -1092 377 -1089 393
rect -1076 377 -1073 393
rect -1060 377 -1057 393
rect -1044 377 -1041 393
rect -652 378 -649 394
rect -613 378 -610 394
rect -584 377 -581 393
rect -568 377 -565 393
rect -552 377 -549 393
rect -536 377 -533 393
rect -308 378 -305 394
rect -269 378 -266 394
rect -240 377 -237 393
rect -224 377 -221 393
rect -208 377 -205 393
rect -192 377 -189 393
rect -50 378 -47 394
rect -11 378 -8 394
rect 18 377 21 393
rect 34 377 37 393
rect 50 377 53 393
rect 66 377 69 393
<< ndiffusion >>
rect -2766 811 -2765 819
rect -2762 811 -2761 819
rect -2696 822 -2694 830
rect -2691 822 -2689 830
rect -2681 822 -2678 830
rect -2675 822 -2672 830
rect -2664 822 -2662 830
rect -2659 822 -2655 830
rect -2647 822 -2645 830
rect -2642 822 -2640 830
rect -2726 810 -2723 818
rect -2720 810 -2718 818
rect -2611 796 -2609 804
rect -2606 796 -2603 804
rect -2595 796 -2593 804
rect -2590 796 -2588 804
rect -2567 796 -2565 804
rect -2562 796 -2560 804
rect -2313 811 -2312 819
rect -2309 811 -2308 819
rect -2243 822 -2241 830
rect -2238 822 -2236 830
rect -2228 822 -2225 830
rect -2222 822 -2219 830
rect -2211 822 -2209 830
rect -2206 822 -2202 830
rect -2194 822 -2192 830
rect -2189 822 -2187 830
rect -2273 810 -2270 818
rect -2267 810 -2265 818
rect -2158 796 -2156 804
rect -2153 796 -2150 804
rect -2142 796 -2140 804
rect -2137 796 -2135 804
rect -2114 796 -2112 804
rect -2109 796 -2107 804
rect -2022 811 -2021 819
rect -2018 811 -2017 819
rect -1952 822 -1950 830
rect -1947 822 -1945 830
rect -1937 822 -1934 830
rect -1931 822 -1928 830
rect -1920 822 -1918 830
rect -1915 822 -1911 830
rect -1903 822 -1901 830
rect -1898 822 -1896 830
rect -1982 810 -1979 818
rect -1976 810 -1974 818
rect -1867 796 -1865 804
rect -1862 796 -1859 804
rect -1851 796 -1849 804
rect -1846 796 -1844 804
rect -1823 796 -1821 804
rect -1818 796 -1816 804
rect -1779 811 -1778 819
rect -1775 811 -1774 819
rect -1709 822 -1707 830
rect -1704 822 -1702 830
rect -1694 822 -1691 830
rect -1688 822 -1685 830
rect -1677 822 -1675 830
rect -1672 822 -1668 830
rect -1660 822 -1658 830
rect -1655 822 -1653 830
rect -1739 810 -1736 818
rect -1733 810 -1731 818
rect -1624 796 -1622 804
rect -1619 796 -1616 804
rect -1608 796 -1606 804
rect -1603 796 -1601 804
rect -1580 796 -1578 804
rect -1575 796 -1573 804
rect -1097 811 -1096 819
rect -1093 811 -1092 819
rect -1027 822 -1025 830
rect -1022 822 -1020 830
rect -1012 822 -1009 830
rect -1006 822 -1003 830
rect -995 822 -993 830
rect -990 822 -986 830
rect -978 822 -976 830
rect -973 822 -971 830
rect -1057 810 -1054 818
rect -1051 810 -1049 818
rect -942 796 -940 804
rect -937 796 -934 804
rect -926 796 -924 804
rect -921 796 -919 804
rect -898 796 -896 804
rect -893 796 -891 804
rect -644 811 -643 819
rect -640 811 -639 819
rect -574 822 -572 830
rect -569 822 -567 830
rect -559 822 -556 830
rect -553 822 -550 830
rect -542 822 -540 830
rect -537 822 -533 830
rect -525 822 -523 830
rect -520 822 -518 830
rect -604 810 -601 818
rect -598 810 -596 818
rect -3090 483 -3087 491
rect -3084 483 -3081 491
rect -3073 483 -3070 491
rect -3067 483 -3064 491
rect -3056 483 -3054 491
rect -3051 483 -3048 491
rect -3040 483 -3038 491
rect -3035 483 -3032 491
rect -3024 483 -3022 491
rect -3019 483 -3017 491
rect -2996 483 -2994 491
rect -2991 483 -2989 491
rect -2962 483 -2959 491
rect -2956 483 -2953 491
rect -2945 483 -2943 491
rect -2940 483 -2937 491
rect -2929 483 -2927 491
rect -2924 483 -2921 491
rect -2913 483 -2911 491
rect -2908 483 -2906 491
rect -2885 483 -2883 491
rect -2880 483 -2878 491
rect -2853 483 -2850 491
rect -2847 483 -2844 491
rect -2836 483 -2834 491
rect -2831 483 -2828 491
rect -2820 483 -2818 491
rect -2815 483 -2813 491
rect -2792 483 -2790 491
rect -2787 483 -2785 491
rect -2754 483 -2751 491
rect -2748 483 -2745 491
rect -2737 483 -2735 491
rect -2732 483 -2730 491
rect -2709 483 -2707 491
rect -2704 483 -2702 491
rect -2675 483 -2673 491
rect -2670 483 -2667 491
rect -2659 483 -2657 491
rect -2654 483 -2651 491
rect -2643 483 -2641 491
rect -2638 483 -2635 491
rect -2627 483 -2625 491
rect -2622 483 -2620 491
rect -2612 483 -2610 491
rect -2607 483 -2605 491
rect -2584 483 -2582 491
rect -2579 483 -2577 491
rect -2519 483 -2516 491
rect -2513 483 -2510 491
rect -2502 483 -2500 491
rect -2497 483 -2494 491
rect -2486 483 -2484 491
rect -2481 483 -2478 491
rect -2470 483 -2468 491
rect -2465 483 -2463 491
rect -2442 483 -2440 491
rect -2437 483 -2435 491
rect -2410 483 -2407 491
rect -2404 483 -2401 491
rect -2393 483 -2391 491
rect -2388 483 -2385 491
rect -2377 483 -2375 491
rect -2372 483 -2370 491
rect -2349 483 -2347 491
rect -2344 483 -2342 491
rect -2311 483 -2308 491
rect -2305 483 -2302 491
rect -2294 483 -2292 491
rect -2289 483 -2287 491
rect -2266 483 -2264 491
rect -2261 483 -2259 491
rect -2232 483 -2230 491
rect -2227 483 -2224 491
rect -2216 483 -2214 491
rect -2211 483 -2208 491
rect -2200 483 -2198 491
rect -2195 483 -2193 491
rect -2185 483 -2182 491
rect -2179 483 -2177 491
rect -2156 483 -2154 491
rect -2151 483 -2149 491
rect -2036 483 -2033 491
rect -2030 483 -2027 491
rect -2019 483 -2017 491
rect -2014 483 -2011 491
rect -2003 483 -2001 491
rect -1998 483 -1996 491
rect -1975 483 -1973 491
rect -1970 483 -1968 491
rect -1937 483 -1934 491
rect -1931 483 -1928 491
rect -1920 483 -1918 491
rect -1915 483 -1913 491
rect -1892 483 -1890 491
rect -1887 483 -1885 491
rect -1835 483 -1833 491
rect -1830 483 -1827 491
rect -1819 483 -1817 491
rect -1814 483 -1811 491
rect -1803 483 -1800 491
rect -1797 483 -1795 491
rect -1774 483 -1772 491
rect -1769 483 -1767 491
rect -1656 481 -1653 489
rect -1650 481 -1647 489
rect -1639 481 -1637 489
rect -1634 481 -1632 489
rect -1611 481 -1609 489
rect -1606 481 -1604 489
rect -1576 481 -1574 489
rect -1571 481 -1568 489
rect -1560 481 -1557 489
rect -1554 481 -1552 489
rect -1531 481 -1529 489
rect -1526 481 -1524 489
rect -2831 274 -2829 282
rect -2826 274 -2824 282
rect -2763 285 -2761 293
rect -2758 285 -2756 293
rect -2748 285 -2745 293
rect -2742 285 -2739 293
rect -2731 285 -2729 293
rect -2726 285 -2723 293
rect -2715 285 -2713 293
rect -2710 285 -2708 293
rect -2793 273 -2790 281
rect -2787 273 -2785 281
rect -489 796 -487 804
rect -484 796 -481 804
rect -473 796 -471 804
rect -468 796 -466 804
rect -445 796 -443 804
rect -440 796 -438 804
rect -353 811 -352 819
rect -349 811 -348 819
rect -283 822 -281 830
rect -278 822 -276 830
rect -268 822 -265 830
rect -262 822 -259 830
rect -251 822 -249 830
rect -246 822 -242 830
rect -234 822 -232 830
rect -229 822 -227 830
rect -313 810 -310 818
rect -307 810 -305 818
rect -198 796 -196 804
rect -193 796 -190 804
rect -182 796 -180 804
rect -177 796 -175 804
rect -154 796 -152 804
rect -149 796 -147 804
rect -110 811 -109 819
rect -106 811 -105 819
rect -40 822 -38 830
rect -35 822 -33 830
rect -25 822 -22 830
rect -19 822 -16 830
rect -8 822 -6 830
rect -3 822 1 830
rect 9 822 11 830
rect 14 822 16 830
rect -70 810 -67 818
rect -64 810 -62 818
rect 45 796 47 804
rect 50 796 53 804
rect 61 796 63 804
rect 66 796 68 804
rect 89 796 91 804
rect 94 796 96 804
rect -1486 481 -1483 489
rect -1480 481 -1477 489
rect -1469 481 -1466 489
rect -1463 481 -1460 489
rect -1452 481 -1450 489
rect -1447 481 -1444 489
rect -1436 481 -1434 489
rect -1431 481 -1428 489
rect -1420 481 -1418 489
rect -1415 481 -1413 489
rect -1392 481 -1390 489
rect -1387 481 -1385 489
rect -1358 481 -1355 489
rect -1352 481 -1349 489
rect -1341 481 -1339 489
rect -1336 481 -1333 489
rect -1325 481 -1323 489
rect -1320 481 -1317 489
rect -1309 481 -1307 489
rect -1304 481 -1302 489
rect -1281 481 -1279 489
rect -1276 481 -1274 489
rect -1249 481 -1246 489
rect -1243 481 -1240 489
rect -1232 481 -1230 489
rect -1227 481 -1224 489
rect -1216 481 -1214 489
rect -1211 481 -1209 489
rect -1188 481 -1186 489
rect -1183 481 -1181 489
rect -1150 481 -1147 489
rect -1144 481 -1141 489
rect -1133 481 -1131 489
rect -1128 481 -1126 489
rect -1105 481 -1103 489
rect -1100 481 -1098 489
rect -1071 481 -1069 489
rect -1066 481 -1063 489
rect -1055 481 -1053 489
rect -1050 481 -1047 489
rect -1039 481 -1037 489
rect -1034 481 -1031 489
rect -1023 481 -1021 489
rect -1018 481 -1016 489
rect -1008 481 -1006 489
rect -1003 481 -1001 489
rect -980 481 -978 489
rect -975 481 -973 489
rect -850 481 -847 489
rect -844 481 -841 489
rect -833 481 -831 489
rect -828 481 -825 489
rect -817 481 -815 489
rect -812 481 -809 489
rect -801 481 -799 489
rect -796 481 -794 489
rect -773 481 -771 489
rect -768 481 -766 489
rect -741 481 -738 489
rect -735 481 -732 489
rect -724 481 -722 489
rect -719 481 -716 489
rect -708 481 -706 489
rect -703 481 -701 489
rect -680 481 -678 489
rect -675 481 -673 489
rect -642 481 -639 489
rect -636 481 -633 489
rect -625 481 -623 489
rect -620 481 -618 489
rect -597 481 -595 489
rect -592 481 -590 489
rect -563 481 -561 489
rect -558 481 -555 489
rect -547 481 -545 489
rect -542 481 -539 489
rect -531 481 -529 489
rect -526 481 -524 489
rect -516 481 -513 489
rect -510 481 -508 489
rect -487 481 -485 489
rect -482 481 -480 489
rect -2323 274 -2321 282
rect -2318 274 -2316 282
rect -2255 285 -2253 293
rect -2250 285 -2248 293
rect -2240 285 -2237 293
rect -2234 285 -2231 293
rect -2223 285 -2221 293
rect -2218 285 -2215 293
rect -2207 285 -2205 293
rect -2202 285 -2200 293
rect -2285 273 -2282 281
rect -2279 273 -2277 281
rect -1979 274 -1977 282
rect -1974 274 -1972 282
rect -1911 285 -1909 293
rect -1906 285 -1904 293
rect -1896 285 -1893 293
rect -1890 285 -1887 293
rect -1879 285 -1877 293
rect -1874 285 -1871 293
rect -1863 285 -1861 293
rect -1858 285 -1856 293
rect -1941 273 -1938 281
rect -1935 273 -1933 281
rect -367 481 -364 489
rect -361 481 -358 489
rect -350 481 -348 489
rect -345 481 -342 489
rect -334 481 -332 489
rect -329 481 -327 489
rect -306 481 -304 489
rect -301 481 -299 489
rect -268 481 -265 489
rect -262 481 -259 489
rect -251 481 -249 489
rect -246 481 -244 489
rect -223 481 -221 489
rect -218 481 -216 489
rect -166 481 -164 489
rect -161 481 -158 489
rect -150 481 -148 489
rect -145 481 -142 489
rect -134 481 -131 489
rect -128 481 -126 489
rect -105 481 -103 489
rect -100 481 -98 489
rect -53 481 -50 489
rect -47 481 -44 489
rect -36 481 -34 489
rect -31 481 -29 489
rect -8 481 -6 489
rect -3 481 -1 489
rect 27 481 29 489
rect 32 481 35 489
rect 43 481 46 489
rect 49 481 51 489
rect 72 481 74 489
rect 77 481 79 489
rect -1598 274 -1596 282
rect -1593 274 -1591 282
rect -1530 285 -1528 293
rect -1525 285 -1523 293
rect -1515 285 -1512 293
rect -1509 285 -1506 293
rect -1498 285 -1496 293
rect -1493 285 -1490 293
rect -1482 285 -1480 293
rect -1477 285 -1475 293
rect -1560 273 -1557 281
rect -1554 273 -1552 281
rect -1162 274 -1160 282
rect -1157 274 -1155 282
rect -1094 285 -1092 293
rect -1089 285 -1087 293
rect -1079 285 -1076 293
rect -1073 285 -1070 293
rect -1062 285 -1060 293
rect -1057 285 -1054 293
rect -1046 285 -1044 293
rect -1041 285 -1037 293
rect -1124 273 -1121 281
rect -1118 273 -1116 281
rect -654 274 -652 282
rect -649 274 -647 282
rect -586 285 -584 293
rect -581 285 -579 293
rect -571 285 -568 293
rect -565 285 -562 293
rect -554 285 -552 293
rect -549 285 -546 293
rect -538 285 -536 293
rect -533 285 -531 293
rect -616 273 -613 281
rect -610 273 -608 281
rect -310 274 -308 282
rect -305 274 -303 282
rect -242 285 -240 293
rect -237 285 -235 293
rect -227 285 -224 293
rect -221 285 -218 293
rect -210 285 -208 293
rect -205 285 -202 293
rect -194 285 -192 293
rect -189 285 -187 293
rect -272 273 -269 281
rect -266 273 -264 281
rect -52 274 -50 282
rect -47 274 -45 282
rect 16 285 18 293
rect 21 285 23 293
rect 31 285 34 293
rect 37 285 40 293
rect 48 285 50 293
rect 53 285 56 293
rect 64 285 66 293
rect 69 285 71 293
rect -14 273 -11 281
rect -8 273 -6 281
<< pdiffusion >>
rect -2766 933 -2765 949
rect -2762 933 -2761 949
rect -2726 933 -2723 949
rect -2720 933 -2718 949
rect -2697 933 -2694 949
rect -2691 933 -2689 949
rect -2681 933 -2678 949
rect -2675 933 -2673 949
rect -2665 933 -2662 949
rect -2659 933 -2656 949
rect -2648 933 -2645 949
rect -2642 933 -2640 949
rect -2610 933 -2609 949
rect -2606 933 -2603 949
rect -2595 933 -2593 949
rect -2590 933 -2588 949
rect -2567 933 -2565 949
rect -2562 933 -2560 949
rect -2313 933 -2312 949
rect -2309 933 -2308 949
rect -2273 933 -2270 949
rect -2267 933 -2265 949
rect -2244 933 -2241 949
rect -2238 933 -2236 949
rect -2228 933 -2225 949
rect -2222 933 -2220 949
rect -2212 933 -2209 949
rect -2206 933 -2203 949
rect -2195 933 -2192 949
rect -2189 933 -2187 949
rect -2157 933 -2156 949
rect -2153 933 -2150 949
rect -2142 933 -2140 949
rect -2137 933 -2135 949
rect -2114 933 -2112 949
rect -2109 933 -2107 949
rect -2022 933 -2021 949
rect -2018 933 -2017 949
rect -1982 933 -1979 949
rect -1976 933 -1974 949
rect -1953 933 -1950 949
rect -1947 933 -1945 949
rect -1937 933 -1934 949
rect -1931 933 -1929 949
rect -1921 933 -1918 949
rect -1915 933 -1912 949
rect -1904 933 -1901 949
rect -1898 933 -1896 949
rect -1866 933 -1865 949
rect -1862 933 -1859 949
rect -1851 933 -1849 949
rect -1846 933 -1844 949
rect -1823 933 -1821 949
rect -1818 933 -1816 949
rect -1779 933 -1778 949
rect -1775 933 -1774 949
rect -1739 933 -1736 949
rect -1733 933 -1731 949
rect -1710 933 -1707 949
rect -1704 933 -1702 949
rect -1694 933 -1691 949
rect -1688 933 -1686 949
rect -1678 933 -1675 949
rect -1672 933 -1669 949
rect -1661 933 -1658 949
rect -1655 933 -1653 949
rect -1623 933 -1622 949
rect -1619 933 -1616 949
rect -1608 933 -1606 949
rect -1603 933 -1601 949
rect -1580 933 -1578 949
rect -1575 933 -1573 949
rect -1097 933 -1096 949
rect -1093 933 -1092 949
rect -1057 933 -1054 949
rect -1051 933 -1049 949
rect -1028 933 -1025 949
rect -1022 933 -1020 949
rect -1012 933 -1009 949
rect -1006 933 -1004 949
rect -996 933 -993 949
rect -990 933 -987 949
rect -979 933 -976 949
rect -973 933 -971 949
rect -941 933 -940 949
rect -937 933 -934 949
rect -926 933 -924 949
rect -921 933 -919 949
rect -898 933 -896 949
rect -893 933 -891 949
rect -644 933 -643 949
rect -640 933 -639 949
rect -604 933 -601 949
rect -598 933 -596 949
rect -575 933 -572 949
rect -569 933 -567 949
rect -559 933 -556 949
rect -553 933 -551 949
rect -543 933 -540 949
rect -537 933 -534 949
rect -526 933 -523 949
rect -520 933 -518 949
rect -488 933 -487 949
rect -484 933 -481 949
rect -473 933 -471 949
rect -468 933 -466 949
rect -445 933 -443 949
rect -440 933 -438 949
rect -353 933 -352 949
rect -349 933 -348 949
rect -313 933 -310 949
rect -307 933 -305 949
rect -284 933 -281 949
rect -278 933 -276 949
rect -268 933 -265 949
rect -262 933 -260 949
rect -252 933 -249 949
rect -246 933 -243 949
rect -235 933 -232 949
rect -229 933 -227 949
rect -197 933 -196 949
rect -193 933 -190 949
rect -182 933 -180 949
rect -177 933 -175 949
rect -154 933 -152 949
rect -149 933 -147 949
rect -110 933 -109 949
rect -106 933 -105 949
rect -70 933 -67 949
rect -64 933 -62 949
rect -41 933 -38 949
rect -35 933 -33 949
rect -25 933 -22 949
rect -19 933 -17 949
rect -9 933 -6 949
rect -3 933 0 949
rect 8 933 11 949
rect 14 933 16 949
rect 46 933 47 949
rect 50 933 53 949
rect 61 933 63 949
rect 66 933 68 949
rect 89 933 91 949
rect 94 933 96 949
rect -3089 601 -3087 617
rect -3084 601 -3080 617
rect -3072 601 -3070 617
rect -3067 601 -3065 617
rect -3057 601 -3054 617
rect -3051 601 -3048 617
rect -3040 601 -3038 617
rect -3035 601 -3032 617
rect -3024 601 -3022 617
rect -3019 601 -3017 617
rect -2996 601 -2994 617
rect -2991 601 -2989 617
rect -2961 601 -2959 617
rect -2956 601 -2954 617
rect -2946 601 -2943 617
rect -2940 601 -2937 617
rect -2929 601 -2927 617
rect -2924 601 -2921 617
rect -2913 601 -2911 617
rect -2908 601 -2906 617
rect -2885 601 -2883 617
rect -2880 601 -2878 617
rect -2852 601 -2850 617
rect -2847 601 -2845 617
rect -2837 601 -2834 617
rect -2831 601 -2828 617
rect -2820 601 -2818 617
rect -2815 601 -2813 617
rect -2792 601 -2790 617
rect -2787 601 -2785 617
rect -2753 601 -2751 617
rect -2748 601 -2745 617
rect -2737 601 -2735 617
rect -2732 601 -2730 617
rect -2709 601 -2707 617
rect -2704 601 -2702 617
rect -2675 601 -2673 617
rect -2670 601 -2667 617
rect -2659 601 -2657 617
rect -2654 601 -2651 617
rect -2643 601 -2641 617
rect -2638 601 -2636 617
rect -2628 601 -2625 617
rect -2622 601 -2621 617
rect -2613 601 -2610 617
rect -2607 601 -2605 617
rect -2584 601 -2582 617
rect -2579 601 -2577 617
rect -2518 601 -2516 617
rect -2513 601 -2511 617
rect -2503 601 -2500 617
rect -2497 601 -2494 617
rect -2486 601 -2484 617
rect -2481 601 -2478 617
rect -2470 601 -2468 617
rect -2465 601 -2463 617
rect -2442 601 -2440 617
rect -2437 601 -2435 617
rect -2409 601 -2407 617
rect -2404 601 -2402 617
rect -2394 601 -2391 617
rect -2388 601 -2385 617
rect -2377 601 -2375 617
rect -2372 601 -2370 617
rect -2349 601 -2347 617
rect -2344 601 -2342 617
rect -2310 601 -2308 617
rect -2305 601 -2302 617
rect -2294 601 -2292 617
rect -2289 601 -2287 617
rect -2266 601 -2264 617
rect -2261 601 -2259 617
rect -2232 601 -2230 617
rect -2227 601 -2224 617
rect -2216 601 -2214 617
rect -2211 601 -2208 617
rect -2200 601 -2198 617
rect -2195 601 -2194 617
rect -2186 601 -2182 617
rect -2179 601 -2177 617
rect -2156 601 -2154 617
rect -2151 601 -2149 617
rect -2035 601 -2033 617
rect -2030 601 -2028 617
rect -2020 601 -2017 617
rect -2014 601 -2011 617
rect -2003 601 -2001 617
rect -1998 601 -1996 617
rect -1975 601 -1973 617
rect -1970 601 -1968 617
rect -1936 601 -1934 617
rect -1931 601 -1928 617
rect -1920 601 -1918 617
rect -1915 601 -1913 617
rect -1892 601 -1890 617
rect -1887 601 -1885 617
rect -1835 601 -1833 617
rect -1830 601 -1827 617
rect -1819 601 -1817 617
rect -1814 601 -1812 617
rect -1804 601 -1800 617
rect -1797 601 -1795 617
rect -1774 601 -1772 617
rect -1769 601 -1767 617
rect -2831 378 -2829 394
rect -2826 378 -2824 394
rect -2793 378 -2790 394
rect -2787 378 -2785 394
rect -1655 599 -1653 615
rect -1650 599 -1647 615
rect -1639 599 -1637 615
rect -1634 599 -1632 615
rect -1611 599 -1609 615
rect -1606 599 -1604 615
rect -1576 599 -1574 615
rect -1571 599 -1569 615
rect -1561 599 -1557 615
rect -1554 599 -1552 615
rect -1531 599 -1529 615
rect -1526 599 -1524 615
rect -1485 599 -1483 615
rect -1480 599 -1476 615
rect -1468 599 -1466 615
rect -1463 599 -1461 615
rect -1453 599 -1450 615
rect -1447 599 -1444 615
rect -1436 599 -1434 615
rect -1431 599 -1428 615
rect -1420 599 -1418 615
rect -1415 599 -1413 615
rect -1392 599 -1390 615
rect -1387 599 -1385 615
rect -1357 599 -1355 615
rect -1352 599 -1350 615
rect -1342 599 -1339 615
rect -1336 599 -1333 615
rect -1325 599 -1323 615
rect -1320 599 -1317 615
rect -1309 599 -1307 615
rect -1304 599 -1302 615
rect -1281 599 -1279 615
rect -1276 599 -1274 615
rect -1248 599 -1246 615
rect -1243 599 -1241 615
rect -1233 599 -1230 615
rect -1227 599 -1224 615
rect -1216 599 -1214 615
rect -1211 599 -1209 615
rect -1188 599 -1186 615
rect -1183 599 -1181 615
rect -1149 599 -1147 615
rect -1144 599 -1141 615
rect -1133 599 -1131 615
rect -1128 599 -1126 615
rect -1105 599 -1103 615
rect -1100 599 -1098 615
rect -1071 599 -1069 615
rect -1066 599 -1063 615
rect -1055 599 -1053 615
rect -1050 599 -1047 615
rect -1039 599 -1037 615
rect -1034 599 -1032 615
rect -1024 599 -1021 615
rect -1018 599 -1017 615
rect -1009 599 -1006 615
rect -1003 599 -1001 615
rect -980 599 -978 615
rect -975 599 -973 615
rect -2764 377 -2761 393
rect -2758 377 -2756 393
rect -2748 377 -2745 393
rect -2742 377 -2740 393
rect -2732 377 -2729 393
rect -2726 377 -2724 393
rect -2716 377 -2713 393
rect -2710 377 -2708 393
rect -2323 378 -2321 394
rect -2318 378 -2316 394
rect -2285 378 -2282 394
rect -2279 378 -2277 394
rect -2256 377 -2253 393
rect -2250 377 -2248 393
rect -2240 377 -2237 393
rect -2234 377 -2232 393
rect -2224 377 -2221 393
rect -2218 377 -2216 393
rect -2208 377 -2205 393
rect -2202 377 -2200 393
rect -1979 378 -1977 394
rect -1974 378 -1972 394
rect -1941 378 -1938 394
rect -1935 378 -1933 394
rect -849 599 -847 615
rect -844 599 -842 615
rect -834 599 -831 615
rect -828 599 -825 615
rect -817 599 -815 615
rect -812 599 -809 615
rect -801 599 -799 615
rect -796 599 -794 615
rect -773 599 -771 615
rect -768 599 -766 615
rect -740 599 -738 615
rect -735 599 -733 615
rect -725 599 -722 615
rect -719 599 -716 615
rect -708 599 -706 615
rect -703 599 -701 615
rect -680 599 -678 615
rect -675 599 -673 615
rect -641 599 -639 615
rect -636 599 -633 615
rect -625 599 -623 615
rect -620 599 -618 615
rect -597 599 -595 615
rect -592 599 -590 615
rect -563 599 -561 615
rect -558 599 -555 615
rect -547 599 -545 615
rect -542 599 -539 615
rect -531 599 -529 615
rect -526 599 -525 615
rect -517 599 -513 615
rect -510 599 -508 615
rect -487 599 -485 615
rect -482 599 -480 615
rect -366 599 -364 615
rect -361 599 -359 615
rect -351 599 -348 615
rect -345 599 -342 615
rect -334 599 -332 615
rect -329 599 -327 615
rect -306 599 -304 615
rect -301 599 -299 615
rect -267 599 -265 615
rect -262 599 -259 615
rect -251 599 -249 615
rect -246 599 -244 615
rect -223 599 -221 615
rect -218 599 -216 615
rect -166 599 -164 615
rect -161 599 -158 615
rect -150 599 -148 615
rect -145 599 -143 615
rect -135 599 -131 615
rect -128 599 -126 615
rect -105 599 -103 615
rect -100 599 -98 615
rect -52 599 -50 615
rect -47 599 -44 615
rect -36 599 -34 615
rect -31 599 -29 615
rect -8 599 -6 615
rect -3 599 -1 615
rect 27 599 29 615
rect 32 599 34 615
rect 42 599 46 615
rect 49 599 51 615
rect 72 599 74 615
rect 77 599 79 615
rect -1912 377 -1909 393
rect -1906 377 -1904 393
rect -1896 377 -1893 393
rect -1890 377 -1888 393
rect -1880 377 -1877 393
rect -1874 377 -1872 393
rect -1864 377 -1861 393
rect -1858 377 -1856 393
rect -1598 378 -1596 394
rect -1593 378 -1591 394
rect -1560 378 -1557 394
rect -1554 378 -1552 394
rect -1531 377 -1528 393
rect -1525 377 -1523 393
rect -1515 377 -1512 393
rect -1509 377 -1507 393
rect -1499 377 -1496 393
rect -1493 377 -1491 393
rect -1483 377 -1480 393
rect -1477 377 -1475 393
rect -1162 378 -1160 394
rect -1157 378 -1155 394
rect -1124 378 -1121 394
rect -1118 378 -1116 394
rect -1095 377 -1092 393
rect -1089 377 -1087 393
rect -1079 377 -1076 393
rect -1073 377 -1071 393
rect -1063 377 -1060 393
rect -1057 377 -1055 393
rect -1047 377 -1044 393
rect -1041 377 -1037 393
rect -654 378 -652 394
rect -649 378 -647 394
rect -616 378 -613 394
rect -610 378 -608 394
rect -587 377 -584 393
rect -581 377 -579 393
rect -571 377 -568 393
rect -565 377 -563 393
rect -555 377 -552 393
rect -549 377 -547 393
rect -539 377 -536 393
rect -533 377 -531 393
rect -310 378 -308 394
rect -305 378 -303 394
rect -272 378 -269 394
rect -266 378 -264 394
rect -243 377 -240 393
rect -237 377 -235 393
rect -227 377 -224 393
rect -221 377 -219 393
rect -211 377 -208 393
rect -205 377 -203 393
rect -195 377 -192 393
rect -189 377 -187 393
rect -52 378 -50 394
rect -47 378 -45 394
rect -14 378 -11 394
rect -8 378 -6 394
rect 15 377 18 393
rect 21 377 23 393
rect 31 377 34 393
rect 37 377 39 393
rect 47 377 50 393
rect 53 377 55 393
rect 63 377 66 393
rect 69 377 71 393
<< ndcontact >>
rect -2774 811 -2766 819
rect -2761 811 -2753 819
rect -2704 822 -2696 830
rect -2689 822 -2681 830
rect -2672 822 -2664 830
rect -2655 822 -2647 830
rect -2640 822 -2632 830
rect -2734 810 -2726 818
rect -2718 810 -2710 818
rect -2619 796 -2611 804
rect -2603 796 -2595 804
rect -2588 796 -2580 804
rect -2575 796 -2567 804
rect -2560 796 -2552 804
rect -2321 811 -2313 819
rect -2308 811 -2300 819
rect -2251 822 -2243 830
rect -2236 822 -2228 830
rect -2219 822 -2211 830
rect -2202 822 -2194 830
rect -2187 822 -2179 830
rect -2281 810 -2273 818
rect -2265 810 -2257 818
rect -2166 796 -2158 804
rect -2150 796 -2142 804
rect -2135 796 -2127 804
rect -2122 796 -2114 804
rect -2107 796 -2099 804
rect -2030 811 -2022 819
rect -2017 811 -2009 819
rect -1960 822 -1952 830
rect -1945 822 -1937 830
rect -1928 822 -1920 830
rect -1911 822 -1903 830
rect -1896 822 -1888 830
rect -1990 810 -1982 818
rect -1974 810 -1966 818
rect -1875 796 -1867 804
rect -1859 796 -1851 804
rect -1844 796 -1836 804
rect -1831 796 -1823 804
rect -1816 796 -1808 804
rect -1787 811 -1779 819
rect -1774 811 -1766 819
rect -1717 822 -1709 830
rect -1702 822 -1694 830
rect -1685 822 -1677 830
rect -1668 822 -1660 830
rect -1653 822 -1645 830
rect -1747 810 -1739 818
rect -1731 810 -1723 818
rect -1632 796 -1624 804
rect -1616 796 -1608 804
rect -1601 796 -1593 804
rect -1588 796 -1580 804
rect -1573 796 -1565 804
rect -1105 811 -1097 819
rect -1092 811 -1084 819
rect -1035 822 -1027 830
rect -1020 822 -1012 830
rect -1003 822 -995 830
rect -986 822 -978 830
rect -971 822 -963 830
rect -1065 810 -1057 818
rect -1049 810 -1041 818
rect -950 796 -942 804
rect -934 796 -926 804
rect -919 796 -911 804
rect -906 796 -898 804
rect -891 796 -883 804
rect -652 811 -644 819
rect -639 811 -631 819
rect -582 822 -574 830
rect -567 822 -559 830
rect -550 822 -542 830
rect -533 822 -525 830
rect -518 822 -510 830
rect -612 810 -604 818
rect -596 810 -588 818
rect -3098 483 -3090 491
rect -3081 483 -3073 491
rect -3064 483 -3056 491
rect -3048 483 -3040 491
rect -3032 483 -3024 491
rect -3017 483 -3009 491
rect -3004 483 -2996 491
rect -2989 483 -2981 491
rect -2970 483 -2962 491
rect -2953 483 -2945 491
rect -2937 483 -2929 491
rect -2921 483 -2913 491
rect -2906 483 -2898 491
rect -2893 483 -2885 491
rect -2878 483 -2870 491
rect -2861 483 -2853 491
rect -2844 483 -2836 491
rect -2828 483 -2820 491
rect -2813 483 -2805 491
rect -2800 483 -2792 491
rect -2785 483 -2777 491
rect -2762 483 -2754 491
rect -2745 483 -2737 491
rect -2730 483 -2722 491
rect -2717 483 -2709 491
rect -2702 483 -2694 491
rect -2683 483 -2675 491
rect -2667 483 -2659 491
rect -2651 483 -2643 491
rect -2635 483 -2627 491
rect -2620 483 -2612 491
rect -2605 483 -2597 491
rect -2592 483 -2584 491
rect -2577 483 -2569 491
rect -2527 483 -2519 491
rect -2510 483 -2502 491
rect -2494 483 -2486 491
rect -2478 483 -2470 491
rect -2463 483 -2455 491
rect -2450 483 -2442 491
rect -2435 483 -2427 491
rect -2418 483 -2410 491
rect -2401 483 -2393 491
rect -2385 483 -2377 491
rect -2370 483 -2362 491
rect -2357 483 -2349 491
rect -2342 483 -2334 491
rect -2319 483 -2311 491
rect -2302 483 -2294 491
rect -2287 483 -2279 491
rect -2274 483 -2266 491
rect -2259 483 -2251 491
rect -2240 483 -2232 491
rect -2224 483 -2216 491
rect -2208 483 -2200 491
rect -2193 483 -2185 491
rect -2177 483 -2169 491
rect -2164 483 -2156 491
rect -2149 483 -2141 491
rect -2044 483 -2036 491
rect -2027 483 -2019 491
rect -2011 483 -2003 491
rect -1996 483 -1988 491
rect -1983 483 -1975 491
rect -1968 483 -1960 491
rect -1945 483 -1937 491
rect -1928 483 -1920 491
rect -1913 483 -1905 491
rect -1900 483 -1892 491
rect -1885 483 -1877 491
rect -1843 483 -1835 491
rect -1827 483 -1819 491
rect -1811 483 -1803 491
rect -1795 483 -1787 491
rect -1782 483 -1774 491
rect -1767 483 -1759 491
rect -1664 481 -1656 489
rect -1647 481 -1639 489
rect -1632 481 -1624 489
rect -1619 481 -1611 489
rect -1604 481 -1596 489
rect -1584 481 -1576 489
rect -1568 481 -1560 489
rect -1552 481 -1544 489
rect -1539 481 -1531 489
rect -1524 481 -1516 489
rect -2839 274 -2831 282
rect -2824 274 -2816 282
rect -2771 285 -2763 293
rect -2756 285 -2748 293
rect -2739 285 -2731 293
rect -2723 285 -2715 293
rect -2708 285 -2700 293
rect -2801 273 -2793 281
rect -2785 273 -2777 281
rect -497 796 -489 804
rect -481 796 -473 804
rect -466 796 -458 804
rect -453 796 -445 804
rect -438 796 -430 804
rect -361 811 -353 819
rect -348 811 -340 819
rect -291 822 -283 830
rect -276 822 -268 830
rect -259 822 -251 830
rect -242 822 -234 830
rect -227 822 -219 830
rect -321 810 -313 818
rect -305 810 -297 818
rect -206 796 -198 804
rect -190 796 -182 804
rect -175 796 -167 804
rect -162 796 -154 804
rect -147 796 -139 804
rect -118 811 -110 819
rect -105 811 -97 819
rect -48 822 -40 830
rect -33 822 -25 830
rect -16 822 -8 830
rect 1 822 9 830
rect 16 822 24 830
rect -78 810 -70 818
rect -62 810 -54 818
rect 37 796 45 804
rect 53 796 61 804
rect 68 796 76 804
rect 81 796 89 804
rect 96 796 104 804
rect -1494 481 -1486 489
rect -1477 481 -1469 489
rect -1460 481 -1452 489
rect -1444 481 -1436 489
rect -1428 481 -1420 489
rect -1413 481 -1405 489
rect -1400 481 -1392 489
rect -1385 481 -1377 489
rect -1366 481 -1358 489
rect -1349 481 -1341 489
rect -1333 481 -1325 489
rect -1317 481 -1309 489
rect -1302 481 -1294 489
rect -1289 481 -1281 489
rect -1274 481 -1266 489
rect -1257 481 -1249 489
rect -1240 481 -1232 489
rect -1224 481 -1216 489
rect -1209 481 -1201 489
rect -1196 481 -1188 489
rect -1181 481 -1173 489
rect -1158 481 -1150 489
rect -1141 481 -1133 489
rect -1126 481 -1118 489
rect -1113 481 -1105 489
rect -1098 481 -1090 489
rect -1079 481 -1071 489
rect -1063 481 -1055 489
rect -1047 481 -1039 489
rect -1031 481 -1023 489
rect -1016 481 -1008 489
rect -1001 481 -993 489
rect -988 481 -980 489
rect -973 481 -965 489
rect -858 481 -850 489
rect -841 481 -833 489
rect -825 481 -817 489
rect -809 481 -801 489
rect -794 481 -786 489
rect -781 481 -773 489
rect -766 481 -758 489
rect -749 481 -741 489
rect -732 481 -724 489
rect -716 481 -708 489
rect -701 481 -693 489
rect -688 481 -680 489
rect -673 481 -665 489
rect -650 481 -642 489
rect -633 481 -625 489
rect -618 481 -610 489
rect -605 481 -597 489
rect -590 481 -582 489
rect -571 481 -563 489
rect -555 481 -547 489
rect -539 481 -531 489
rect -524 481 -516 489
rect -508 481 -500 489
rect -495 481 -487 489
rect -480 481 -472 489
rect -2331 274 -2323 282
rect -2316 274 -2308 282
rect -2263 285 -2255 293
rect -2248 285 -2240 293
rect -2231 285 -2223 293
rect -2215 285 -2207 293
rect -2200 285 -2192 293
rect -2293 273 -2285 281
rect -2277 273 -2269 281
rect -1987 274 -1979 282
rect -1972 274 -1964 282
rect -1919 285 -1911 293
rect -1904 285 -1896 293
rect -1887 285 -1879 293
rect -1871 285 -1863 293
rect -1856 285 -1848 293
rect -1949 273 -1941 281
rect -1933 273 -1925 281
rect -375 481 -367 489
rect -358 481 -350 489
rect -342 481 -334 489
rect -327 481 -319 489
rect -314 481 -306 489
rect -299 481 -291 489
rect -276 481 -268 489
rect -259 481 -251 489
rect -244 481 -236 489
rect -231 481 -223 489
rect -216 481 -208 489
rect -174 481 -166 489
rect -158 481 -150 489
rect -142 481 -134 489
rect -126 481 -118 489
rect -113 481 -105 489
rect -98 481 -90 489
rect -61 481 -53 489
rect -44 481 -36 489
rect -29 481 -21 489
rect -16 481 -8 489
rect -1 481 7 489
rect 19 481 27 489
rect 35 481 43 489
rect 51 481 59 489
rect 64 481 72 489
rect 79 481 87 489
rect -1606 274 -1598 282
rect -1591 274 -1583 282
rect -1538 285 -1530 293
rect -1523 285 -1515 293
rect -1506 285 -1498 293
rect -1490 285 -1482 293
rect -1475 285 -1467 293
rect -1568 273 -1560 281
rect -1552 273 -1544 281
rect -1170 274 -1162 282
rect -1155 274 -1147 282
rect -1102 285 -1094 293
rect -1087 285 -1079 293
rect -1070 285 -1062 293
rect -1054 285 -1046 293
rect -1037 285 -1029 293
rect -1132 273 -1124 281
rect -1116 273 -1108 281
rect -662 274 -654 282
rect -647 274 -639 282
rect -594 285 -586 293
rect -579 285 -571 293
rect -562 285 -554 293
rect -546 285 -538 293
rect -531 285 -523 293
rect -624 273 -616 281
rect -608 273 -600 281
rect -318 274 -310 282
rect -303 274 -295 282
rect -250 285 -242 293
rect -235 285 -227 293
rect -218 285 -210 293
rect -202 285 -194 293
rect -187 285 -179 293
rect -280 273 -272 281
rect -264 273 -256 281
rect -60 274 -52 282
rect -45 274 -37 282
rect 8 285 16 293
rect 23 285 31 293
rect 40 285 48 293
rect 56 285 64 293
rect 71 285 79 293
rect -22 273 -14 281
rect -6 273 2 281
<< pdcontact >>
rect -2774 933 -2766 949
rect -2761 933 -2753 949
rect -2734 933 -2726 949
rect -2718 933 -2710 949
rect -2705 933 -2697 949
rect -2689 933 -2681 949
rect -2673 933 -2665 949
rect -2656 933 -2648 949
rect -2640 933 -2632 949
rect -2618 933 -2610 949
rect -2603 933 -2595 949
rect -2588 933 -2580 949
rect -2575 933 -2567 949
rect -2560 933 -2552 949
rect -2321 933 -2313 949
rect -2308 933 -2300 949
rect -2281 933 -2273 949
rect -2265 933 -2257 949
rect -2252 933 -2244 949
rect -2236 933 -2228 949
rect -2220 933 -2212 949
rect -2203 933 -2195 949
rect -2187 933 -2179 949
rect -2165 933 -2157 949
rect -2150 933 -2142 949
rect -2135 933 -2127 949
rect -2122 933 -2114 949
rect -2107 933 -2099 949
rect -2030 933 -2022 949
rect -2017 933 -2009 949
rect -1990 933 -1982 949
rect -1974 933 -1966 949
rect -1961 933 -1953 949
rect -1945 933 -1937 949
rect -1929 933 -1921 949
rect -1912 933 -1904 949
rect -1896 933 -1888 949
rect -1874 933 -1866 949
rect -1859 933 -1851 949
rect -1844 933 -1836 949
rect -1831 933 -1823 949
rect -1816 933 -1808 949
rect -1787 933 -1779 949
rect -1774 933 -1766 949
rect -1747 933 -1739 949
rect -1731 933 -1723 949
rect -1718 933 -1710 949
rect -1702 933 -1694 949
rect -1686 933 -1678 949
rect -1669 933 -1661 949
rect -1653 933 -1645 949
rect -1631 933 -1623 949
rect -1616 933 -1608 949
rect -1601 933 -1593 949
rect -1588 933 -1580 949
rect -1573 933 -1565 949
rect -1105 933 -1097 949
rect -1092 933 -1084 949
rect -1065 933 -1057 949
rect -1049 933 -1041 949
rect -1036 933 -1028 949
rect -1020 933 -1012 949
rect -1004 933 -996 949
rect -987 933 -979 949
rect -971 933 -963 949
rect -949 933 -941 949
rect -934 933 -926 949
rect -919 933 -911 949
rect -906 933 -898 949
rect -891 933 -883 949
rect -652 933 -644 949
rect -639 933 -631 949
rect -612 933 -604 949
rect -596 933 -588 949
rect -583 933 -575 949
rect -567 933 -559 949
rect -551 933 -543 949
rect -534 933 -526 949
rect -518 933 -510 949
rect -496 933 -488 949
rect -481 933 -473 949
rect -466 933 -458 949
rect -453 933 -445 949
rect -438 933 -430 949
rect -361 933 -353 949
rect -348 933 -340 949
rect -321 933 -313 949
rect -305 933 -297 949
rect -292 933 -284 949
rect -276 933 -268 949
rect -260 933 -252 949
rect -243 933 -235 949
rect -227 933 -219 949
rect -205 933 -197 949
rect -190 933 -182 949
rect -175 933 -167 949
rect -162 933 -154 949
rect -147 933 -139 949
rect -118 933 -110 949
rect -105 933 -97 949
rect -78 933 -70 949
rect -62 933 -54 949
rect -49 933 -41 949
rect -33 933 -25 949
rect -17 933 -9 949
rect 0 933 8 949
rect 16 933 24 949
rect 38 933 46 949
rect 53 933 61 949
rect 68 933 76 949
rect 81 933 89 949
rect 96 933 104 949
rect -3097 601 -3089 617
rect -3080 601 -3072 617
rect -3065 601 -3057 617
rect -3048 601 -3040 617
rect -3032 601 -3024 617
rect -3017 601 -3009 617
rect -3004 601 -2996 617
rect -2989 601 -2981 617
rect -2969 601 -2961 617
rect -2954 601 -2946 617
rect -2937 601 -2929 617
rect -2921 601 -2913 617
rect -2906 601 -2898 617
rect -2893 601 -2885 617
rect -2878 601 -2870 617
rect -2860 601 -2852 617
rect -2845 601 -2837 617
rect -2828 601 -2820 617
rect -2813 601 -2805 617
rect -2800 601 -2792 617
rect -2785 601 -2777 617
rect -2761 601 -2753 617
rect -2745 601 -2737 617
rect -2730 601 -2722 617
rect -2717 601 -2709 617
rect -2702 601 -2694 617
rect -2683 601 -2675 617
rect -2667 601 -2659 617
rect -2651 601 -2643 617
rect -2636 601 -2628 617
rect -2621 601 -2613 617
rect -2605 601 -2597 617
rect -2592 601 -2584 617
rect -2577 601 -2569 617
rect -2526 601 -2518 617
rect -2511 601 -2503 617
rect -2494 601 -2486 617
rect -2478 601 -2470 617
rect -2463 601 -2455 617
rect -2450 601 -2442 617
rect -2435 601 -2427 617
rect -2417 601 -2409 617
rect -2402 601 -2394 617
rect -2385 601 -2377 617
rect -2370 601 -2362 617
rect -2357 601 -2349 617
rect -2342 601 -2334 617
rect -2318 601 -2310 617
rect -2302 601 -2294 617
rect -2287 601 -2279 617
rect -2274 601 -2266 617
rect -2259 601 -2251 617
rect -2240 601 -2232 617
rect -2224 601 -2216 617
rect -2208 601 -2200 617
rect -2194 601 -2186 617
rect -2177 601 -2169 617
rect -2164 601 -2156 617
rect -2149 601 -2141 617
rect -2043 601 -2035 617
rect -2028 601 -2020 617
rect -2011 601 -2003 617
rect -1996 601 -1988 617
rect -1983 601 -1975 617
rect -1968 601 -1960 617
rect -1944 601 -1936 617
rect -1928 601 -1920 617
rect -1913 601 -1905 617
rect -1900 601 -1892 617
rect -1885 601 -1877 617
rect -1843 601 -1835 617
rect -1827 601 -1819 617
rect -1812 601 -1804 617
rect -1795 601 -1787 617
rect -1782 601 -1774 617
rect -1767 601 -1759 617
rect -2839 378 -2831 394
rect -2824 378 -2816 394
rect -2801 378 -2793 394
rect -2785 378 -2777 394
rect -1663 599 -1655 615
rect -1647 599 -1639 615
rect -1632 599 -1624 615
rect -1619 599 -1611 615
rect -1604 599 -1596 615
rect -1584 599 -1576 615
rect -1569 599 -1561 615
rect -1552 599 -1544 615
rect -1539 599 -1531 615
rect -1524 599 -1516 615
rect -1493 599 -1485 615
rect -1476 599 -1468 615
rect -1461 599 -1453 615
rect -1444 599 -1436 615
rect -1428 599 -1420 615
rect -1413 599 -1405 615
rect -1400 599 -1392 615
rect -1385 599 -1377 615
rect -1365 599 -1357 615
rect -1350 599 -1342 615
rect -1333 599 -1325 615
rect -1317 599 -1309 615
rect -1302 599 -1294 615
rect -1289 599 -1281 615
rect -1274 599 -1266 615
rect -1256 599 -1248 615
rect -1241 599 -1233 615
rect -1224 599 -1216 615
rect -1209 599 -1201 615
rect -1196 599 -1188 615
rect -1181 599 -1173 615
rect -1157 599 -1149 615
rect -1141 599 -1133 615
rect -1126 599 -1118 615
rect -1113 599 -1105 615
rect -1098 599 -1090 615
rect -1079 599 -1071 615
rect -1063 599 -1055 615
rect -1047 599 -1039 615
rect -1032 599 -1024 615
rect -1017 599 -1009 615
rect -1001 599 -993 615
rect -988 599 -980 615
rect -973 599 -965 615
rect -2772 377 -2764 393
rect -2756 377 -2748 393
rect -2740 377 -2732 393
rect -2724 377 -2716 393
rect -2708 377 -2700 393
rect -2331 378 -2323 394
rect -2316 378 -2308 394
rect -2293 378 -2285 394
rect -2277 378 -2269 394
rect -2264 377 -2256 393
rect -2248 377 -2240 393
rect -2232 377 -2224 393
rect -2216 377 -2208 393
rect -2200 377 -2192 393
rect -1987 378 -1979 394
rect -1972 378 -1964 394
rect -1949 378 -1941 394
rect -1933 378 -1925 394
rect -857 599 -849 615
rect -842 599 -834 615
rect -825 599 -817 615
rect -809 599 -801 615
rect -794 599 -786 615
rect -781 599 -773 615
rect -766 599 -758 615
rect -748 599 -740 615
rect -733 599 -725 615
rect -716 599 -708 615
rect -701 599 -693 615
rect -688 599 -680 615
rect -673 599 -665 615
rect -649 599 -641 615
rect -633 599 -625 615
rect -618 599 -610 615
rect -605 599 -597 615
rect -590 599 -582 615
rect -571 599 -563 615
rect -555 599 -547 615
rect -539 599 -531 615
rect -525 599 -517 615
rect -508 599 -500 615
rect -495 599 -487 615
rect -480 599 -472 615
rect -374 599 -366 615
rect -359 599 -351 615
rect -342 599 -334 615
rect -327 599 -319 615
rect -314 599 -306 615
rect -299 599 -291 615
rect -275 599 -267 615
rect -259 599 -251 615
rect -244 599 -236 615
rect -231 599 -223 615
rect -216 599 -208 615
rect -174 599 -166 615
rect -158 599 -150 615
rect -143 599 -135 615
rect -126 599 -118 615
rect -113 599 -105 615
rect -98 599 -90 615
rect -60 599 -52 615
rect -44 599 -36 615
rect -29 599 -21 615
rect -16 599 -8 615
rect -1 599 7 615
rect 19 599 27 615
rect 34 599 42 615
rect 51 599 59 615
rect 64 599 72 615
rect 79 599 87 615
rect -1920 377 -1912 393
rect -1904 377 -1896 393
rect -1888 377 -1880 393
rect -1872 377 -1864 393
rect -1856 377 -1848 393
rect -1606 378 -1598 394
rect -1591 378 -1583 394
rect -1568 378 -1560 394
rect -1552 378 -1544 394
rect -1539 377 -1531 393
rect -1523 377 -1515 393
rect -1507 377 -1499 393
rect -1491 377 -1483 393
rect -1475 377 -1467 393
rect -1170 378 -1162 394
rect -1155 378 -1147 394
rect -1132 378 -1124 394
rect -1116 378 -1108 394
rect -1103 377 -1095 393
rect -1087 377 -1079 393
rect -1071 377 -1063 393
rect -1055 377 -1047 393
rect -1037 377 -1029 393
rect -662 378 -654 394
rect -647 378 -639 394
rect -624 378 -616 394
rect -608 378 -600 394
rect -595 377 -587 393
rect -579 377 -571 393
rect -563 377 -555 393
rect -547 377 -539 393
rect -531 377 -523 393
rect -318 378 -310 394
rect -303 378 -295 394
rect -280 378 -272 394
rect -264 378 -256 394
rect -251 377 -243 393
rect -235 377 -227 393
rect -219 377 -211 393
rect -203 377 -195 393
rect -187 377 -179 393
rect -60 378 -52 394
rect -45 378 -37 394
rect -22 378 -14 394
rect -6 378 2 394
rect 7 377 15 393
rect 23 377 31 393
rect 39 377 47 393
rect 55 377 63 393
rect 71 377 79 393
<< psubstratepcontact >>
rect -2774 783 -2766 791
rect -2760 783 -2752 791
rect -2734 783 -2726 791
rect -2717 783 -2709 791
rect -2704 783 -2696 791
rect -2687 783 -2679 791
rect -2655 783 -2647 791
rect -2638 783 -2630 791
rect -2619 783 -2611 791
rect -2603 783 -2595 791
rect -2588 783 -2580 791
rect -2575 783 -2567 791
rect -2560 783 -2552 791
rect -2321 783 -2313 791
rect -2307 783 -2299 791
rect -2281 783 -2273 791
rect -2264 783 -2256 791
rect -2251 783 -2243 791
rect -2234 783 -2226 791
rect -2202 783 -2194 791
rect -2185 783 -2177 791
rect -2166 783 -2158 791
rect -2150 783 -2142 791
rect -2135 783 -2127 791
rect -2122 783 -2114 791
rect -2107 783 -2099 791
rect -2030 783 -2022 791
rect -2016 783 -2008 791
rect -1990 783 -1982 791
rect -1973 783 -1965 791
rect -1960 783 -1952 791
rect -1943 783 -1935 791
rect -1911 783 -1903 791
rect -1894 783 -1886 791
rect -1875 783 -1867 791
rect -1859 783 -1851 791
rect -1844 783 -1836 791
rect -1831 783 -1823 791
rect -1816 783 -1808 791
rect -1787 783 -1779 791
rect -1773 783 -1765 791
rect -1747 783 -1739 791
rect -1730 783 -1722 791
rect -1717 783 -1709 791
rect -1700 783 -1692 791
rect -1668 783 -1660 791
rect -1651 783 -1643 791
rect -1632 783 -1624 791
rect -1616 783 -1608 791
rect -1601 783 -1593 791
rect -1588 783 -1580 791
rect -1573 783 -1565 791
rect -1105 783 -1097 791
rect -1091 783 -1083 791
rect -1065 783 -1057 791
rect -1048 783 -1040 791
rect -1035 783 -1027 791
rect -1018 783 -1010 791
rect -986 783 -978 791
rect -969 783 -961 791
rect -950 783 -942 791
rect -934 783 -926 791
rect -919 783 -911 791
rect -906 783 -898 791
rect -891 783 -883 791
rect -652 783 -644 791
rect -638 783 -630 791
rect -612 783 -604 791
rect -595 783 -587 791
rect -582 783 -574 791
rect -565 783 -557 791
rect -533 783 -525 791
rect -516 783 -508 791
rect -3098 470 -3090 478
rect -3081 470 -3073 478
rect -3064 470 -3056 478
rect -3048 470 -3040 478
rect -3032 470 -3024 478
rect -3017 470 -3009 478
rect -3004 470 -2996 478
rect -2989 470 -2981 478
rect -2970 470 -2962 478
rect -2953 470 -2945 478
rect -2937 470 -2929 478
rect -2921 470 -2913 478
rect -2906 470 -2898 478
rect -2893 470 -2885 478
rect -2878 470 -2870 478
rect -2861 470 -2853 478
rect -2844 470 -2836 478
rect -2828 470 -2820 478
rect -2813 470 -2805 478
rect -2800 470 -2792 478
rect -2785 470 -2777 478
rect -2762 470 -2754 478
rect -2745 470 -2737 478
rect -2730 470 -2722 478
rect -2717 470 -2709 478
rect -2702 470 -2694 478
rect -2683 470 -2675 478
rect -2667 470 -2659 478
rect -2651 470 -2643 478
rect -2635 470 -2627 478
rect -2620 470 -2612 478
rect -2605 470 -2597 478
rect -2592 470 -2584 478
rect -2577 470 -2569 478
rect -2527 470 -2519 478
rect -2510 470 -2502 478
rect -2494 470 -2486 478
rect -2478 470 -2470 478
rect -2463 470 -2455 478
rect -2450 470 -2442 478
rect -2435 470 -2427 478
rect -2418 470 -2410 478
rect -2401 470 -2393 478
rect -2385 470 -2377 478
rect -2370 470 -2362 478
rect -2357 470 -2349 478
rect -2342 470 -2334 478
rect -2319 470 -2311 478
rect -2302 470 -2294 478
rect -2287 470 -2279 478
rect -2274 470 -2266 478
rect -2259 470 -2251 478
rect -2240 470 -2232 478
rect -2224 470 -2216 478
rect -2208 470 -2200 478
rect -2193 470 -2185 478
rect -2177 470 -2169 478
rect -2164 470 -2156 478
rect -2149 470 -2141 478
rect -2044 470 -2036 478
rect -2027 470 -2019 478
rect -2011 470 -2003 478
rect -1996 470 -1988 478
rect -1983 470 -1975 478
rect -1968 470 -1960 478
rect -1945 470 -1937 478
rect -1928 470 -1920 478
rect -1913 470 -1905 478
rect -1900 470 -1892 478
rect -1885 470 -1877 478
rect -1843 470 -1835 478
rect -1827 470 -1819 478
rect -1811 470 -1803 478
rect -1795 470 -1787 478
rect -1782 470 -1774 478
rect -1767 470 -1759 478
rect -1664 468 -1656 476
rect -1647 468 -1639 476
rect -1632 468 -1624 476
rect -1619 468 -1611 476
rect -1604 468 -1596 476
rect -1584 468 -1576 476
rect -1568 468 -1560 476
rect -1552 468 -1544 476
rect -1539 468 -1531 476
rect -1524 468 -1516 476
rect -497 783 -489 791
rect -481 783 -473 791
rect -466 783 -458 791
rect -453 783 -445 791
rect -438 783 -430 791
rect -361 783 -353 791
rect -347 783 -339 791
rect -321 783 -313 791
rect -304 783 -296 791
rect -291 783 -283 791
rect -274 783 -266 791
rect -242 783 -234 791
rect -225 783 -217 791
rect -206 783 -198 791
rect -190 783 -182 791
rect -175 783 -167 791
rect -162 783 -154 791
rect -147 783 -139 791
rect -118 783 -110 791
rect -104 783 -96 791
rect -78 783 -70 791
rect -61 783 -53 791
rect -48 783 -40 791
rect -31 783 -23 791
rect 1 783 9 791
rect 18 783 26 791
rect 37 783 45 791
rect 53 783 61 791
rect 68 783 76 791
rect 81 783 89 791
rect 96 783 104 791
rect -1494 468 -1486 476
rect -1477 468 -1469 476
rect -1460 468 -1452 476
rect -1444 468 -1436 476
rect -1428 468 -1420 476
rect -1413 468 -1405 476
rect -1400 468 -1392 476
rect -1385 468 -1377 476
rect -1366 468 -1358 476
rect -1349 468 -1341 476
rect -1333 468 -1325 476
rect -1317 468 -1309 476
rect -1302 468 -1294 476
rect -1289 468 -1281 476
rect -1274 468 -1266 476
rect -1257 468 -1249 476
rect -1240 468 -1232 476
rect -1224 468 -1216 476
rect -1209 468 -1201 476
rect -1196 468 -1188 476
rect -1181 468 -1173 476
rect -1158 468 -1150 476
rect -1141 468 -1133 476
rect -1126 468 -1118 476
rect -1113 468 -1105 476
rect -1098 468 -1090 476
rect -1079 468 -1071 476
rect -1063 468 -1055 476
rect -1047 468 -1039 476
rect -1031 468 -1023 476
rect -1016 468 -1008 476
rect -1001 468 -993 476
rect -988 468 -980 476
rect -973 468 -965 476
rect -858 468 -850 476
rect -841 468 -833 476
rect -825 468 -817 476
rect -809 468 -801 476
rect -794 468 -786 476
rect -781 468 -773 476
rect -766 468 -758 476
rect -749 468 -741 476
rect -732 468 -724 476
rect -716 468 -708 476
rect -701 468 -693 476
rect -688 468 -680 476
rect -673 468 -665 476
rect -650 468 -642 476
rect -633 468 -625 476
rect -618 468 -610 476
rect -605 468 -597 476
rect -590 468 -582 476
rect -571 468 -563 476
rect -555 468 -547 476
rect -539 468 -531 476
rect -524 468 -516 476
rect -508 468 -500 476
rect -495 468 -487 476
rect -480 468 -472 476
rect -375 468 -367 476
rect -358 468 -350 476
rect -342 468 -334 476
rect -327 468 -319 476
rect -314 468 -306 476
rect -299 468 -291 476
rect -276 468 -268 476
rect -259 468 -251 476
rect -244 468 -236 476
rect -231 468 -223 476
rect -216 468 -208 476
rect -174 468 -166 476
rect -158 468 -150 476
rect -142 468 -134 476
rect -126 468 -118 476
rect -113 468 -105 476
rect -98 468 -90 476
rect -61 468 -53 476
rect -44 468 -36 476
rect -29 468 -21 476
rect -16 468 -8 476
rect -1 468 7 476
rect 19 468 27 476
rect 35 468 43 476
rect 51 468 59 476
rect 64 468 72 476
rect 79 468 87 476
rect -2839 246 -2831 254
rect -2823 246 -2815 254
rect -2801 246 -2793 254
rect -2784 246 -2776 254
rect -2771 246 -2763 254
rect -2754 246 -2746 254
rect -2723 246 -2715 254
rect -2706 246 -2698 254
rect -2331 246 -2323 254
rect -2315 246 -2307 254
rect -2293 246 -2285 254
rect -2276 246 -2268 254
rect -2263 246 -2255 254
rect -2246 246 -2238 254
rect -2215 246 -2207 254
rect -2198 246 -2190 254
rect -1987 246 -1979 254
rect -1971 246 -1963 254
rect -1949 246 -1941 254
rect -1932 246 -1924 254
rect -1919 246 -1911 254
rect -1902 246 -1894 254
rect -1871 246 -1863 254
rect -1854 246 -1846 254
rect -1606 246 -1598 254
rect -1590 246 -1582 254
rect -1568 246 -1560 254
rect -1551 246 -1543 254
rect -1538 246 -1530 254
rect -1521 246 -1513 254
rect -1490 246 -1482 254
rect -1473 246 -1465 254
rect -1170 246 -1162 254
rect -1154 246 -1146 254
rect -1132 246 -1124 254
rect -1115 246 -1107 254
rect -1102 246 -1094 254
rect -1085 246 -1077 254
rect -1054 246 -1046 254
rect -1037 246 -1029 254
rect -662 246 -654 254
rect -646 246 -638 254
rect -624 246 -616 254
rect -607 246 -599 254
rect -594 246 -586 254
rect -577 246 -569 254
rect -546 246 -538 254
rect -529 246 -521 254
rect -318 246 -310 254
rect -302 246 -294 254
rect -280 246 -272 254
rect -263 246 -255 254
rect -250 246 -242 254
rect -233 246 -225 254
rect -202 246 -194 254
rect -185 246 -177 254
rect -60 246 -52 254
rect -44 246 -36 254
rect -22 246 -14 254
rect -5 246 3 254
rect 8 246 16 254
rect 25 246 33 254
rect 56 246 64 254
rect 73 246 81 254
<< nsubstratencontact >>
rect -2774 957 -2766 965
rect -2761 957 -2753 965
rect -2734 957 -2726 965
rect -2718 957 -2710 965
rect -2705 957 -2697 965
rect -2689 957 -2681 965
rect -2656 957 -2648 965
rect -2640 957 -2632 965
rect -2618 957 -2610 965
rect -2603 957 -2595 965
rect -2588 957 -2580 965
rect -2575 957 -2567 965
rect -2560 957 -2552 965
rect -2321 957 -2313 965
rect -2308 957 -2300 965
rect -2281 957 -2273 965
rect -2265 957 -2257 965
rect -2252 957 -2244 965
rect -2236 957 -2228 965
rect -2203 957 -2195 965
rect -2187 957 -2179 965
rect -2165 957 -2157 965
rect -2150 957 -2142 965
rect -2135 957 -2127 965
rect -2122 957 -2114 965
rect -2107 957 -2099 965
rect -2030 957 -2022 965
rect -2017 957 -2009 965
rect -1990 957 -1982 965
rect -1974 957 -1966 965
rect -1961 957 -1953 965
rect -1945 957 -1937 965
rect -1912 957 -1904 965
rect -1896 957 -1888 965
rect -1874 957 -1866 965
rect -1859 957 -1851 965
rect -1844 957 -1836 965
rect -1831 957 -1823 965
rect -1816 957 -1808 965
rect -1787 957 -1779 965
rect -1774 957 -1766 965
rect -1747 957 -1739 965
rect -1731 957 -1723 965
rect -1718 957 -1710 965
rect -1702 957 -1694 965
rect -1669 957 -1661 965
rect -1653 957 -1645 965
rect -1631 957 -1623 965
rect -1616 957 -1608 965
rect -1601 957 -1593 965
rect -1588 957 -1580 965
rect -1573 957 -1565 965
rect -1105 957 -1097 965
rect -1092 957 -1084 965
rect -1065 957 -1057 965
rect -1049 957 -1041 965
rect -1036 957 -1028 965
rect -1020 957 -1012 965
rect -987 957 -979 965
rect -971 957 -963 965
rect -949 957 -941 965
rect -934 957 -926 965
rect -919 957 -911 965
rect -906 957 -898 965
rect -891 957 -883 965
rect -652 957 -644 965
rect -639 957 -631 965
rect -612 957 -604 965
rect -596 957 -588 965
rect -583 957 -575 965
rect -567 957 -559 965
rect -534 957 -526 965
rect -518 957 -510 965
rect -496 957 -488 965
rect -481 957 -473 965
rect -466 957 -458 965
rect -453 957 -445 965
rect -438 957 -430 965
rect -361 957 -353 965
rect -348 957 -340 965
rect -321 957 -313 965
rect -305 957 -297 965
rect -292 957 -284 965
rect -276 957 -268 965
rect -243 957 -235 965
rect -227 957 -219 965
rect -205 957 -197 965
rect -190 957 -182 965
rect -175 957 -167 965
rect -162 957 -154 965
rect -147 957 -139 965
rect -118 957 -110 965
rect -105 957 -97 965
rect -78 957 -70 965
rect -62 957 -54 965
rect -49 957 -41 965
rect -33 957 -25 965
rect 0 957 8 965
rect 16 957 24 965
rect 38 957 46 965
rect 53 957 61 965
rect 68 957 76 965
rect 81 957 89 965
rect 96 957 104 965
rect -3097 625 -3089 633
rect -3080 625 -3072 633
rect -3065 625 -3057 633
rect -3048 625 -3040 633
rect -3032 625 -3024 633
rect -3017 625 -3009 633
rect -3004 625 -2996 633
rect -2989 625 -2981 633
rect -2969 625 -2961 633
rect -2954 625 -2946 633
rect -2937 625 -2929 633
rect -2921 625 -2913 633
rect -2906 625 -2898 633
rect -2893 625 -2885 633
rect -2878 625 -2870 633
rect -2860 625 -2852 633
rect -2845 625 -2837 633
rect -2828 625 -2820 633
rect -2813 625 -2805 633
rect -2800 625 -2792 633
rect -2785 625 -2777 633
rect -2761 625 -2753 633
rect -2745 625 -2737 633
rect -2730 625 -2722 633
rect -2717 625 -2709 633
rect -2702 625 -2694 633
rect -2683 625 -2675 633
rect -2667 625 -2659 633
rect -2636 625 -2628 633
rect -2621 625 -2613 633
rect -2605 625 -2597 633
rect -2592 625 -2584 633
rect -2577 625 -2569 633
rect -2526 625 -2518 633
rect -2511 625 -2503 633
rect -2494 625 -2486 633
rect -2478 625 -2470 633
rect -2463 625 -2455 633
rect -2450 625 -2442 633
rect -2435 625 -2427 633
rect -2417 625 -2409 633
rect -2402 625 -2394 633
rect -2385 625 -2377 633
rect -2370 625 -2362 633
rect -2357 625 -2349 633
rect -2342 625 -2334 633
rect -2318 625 -2310 633
rect -2302 625 -2294 633
rect -2287 625 -2279 633
rect -2274 625 -2266 633
rect -2259 625 -2251 633
rect -2240 625 -2232 633
rect -2224 625 -2216 633
rect -2194 625 -2186 633
rect -2177 625 -2169 633
rect -2164 625 -2156 633
rect -2149 625 -2141 633
rect -2043 625 -2035 633
rect -2028 625 -2020 633
rect -2011 625 -2003 633
rect -1996 625 -1988 633
rect -1983 625 -1975 633
rect -1968 625 -1960 633
rect -1944 625 -1936 633
rect -1928 625 -1920 633
rect -1913 625 -1905 633
rect -1900 625 -1892 633
rect -1885 625 -1877 633
rect -1843 625 -1835 633
rect -1827 625 -1819 633
rect -1812 625 -1804 633
rect -1795 625 -1787 633
rect -1782 625 -1774 633
rect -1767 625 -1759 633
rect -1663 623 -1655 631
rect -1647 623 -1639 631
rect -1632 623 -1624 631
rect -1619 623 -1611 631
rect -1604 623 -1596 631
rect -1584 623 -1576 631
rect -1569 623 -1561 631
rect -1552 623 -1544 631
rect -1539 623 -1531 631
rect -1524 623 -1516 631
rect -1493 623 -1485 631
rect -1476 623 -1468 631
rect -1461 623 -1453 631
rect -1444 623 -1436 631
rect -1428 623 -1420 631
rect -1413 623 -1405 631
rect -1400 623 -1392 631
rect -1385 623 -1377 631
rect -1365 623 -1357 631
rect -1350 623 -1342 631
rect -1333 623 -1325 631
rect -1317 623 -1309 631
rect -1302 623 -1294 631
rect -1289 623 -1281 631
rect -1274 623 -1266 631
rect -1256 623 -1248 631
rect -1241 623 -1233 631
rect -1224 623 -1216 631
rect -1209 623 -1201 631
rect -1196 623 -1188 631
rect -1181 623 -1173 631
rect -1157 623 -1149 631
rect -1141 623 -1133 631
rect -1126 623 -1118 631
rect -1113 623 -1105 631
rect -1098 623 -1090 631
rect -1079 623 -1071 631
rect -1063 623 -1055 631
rect -1032 623 -1024 631
rect -1017 623 -1009 631
rect -1001 623 -993 631
rect -988 623 -980 631
rect -973 623 -965 631
rect -2839 402 -2831 410
rect -2824 402 -2816 410
rect -2801 402 -2793 410
rect -2785 402 -2777 410
rect -2772 402 -2764 410
rect -2756 402 -2748 410
rect -2724 402 -2716 410
rect -2708 402 -2700 410
rect -2331 402 -2323 410
rect -2316 402 -2308 410
rect -2293 402 -2285 410
rect -2277 402 -2269 410
rect -2264 402 -2256 410
rect -2248 402 -2240 410
rect -2216 402 -2208 410
rect -2200 402 -2192 410
rect -1987 402 -1979 410
rect -1972 402 -1964 410
rect -1949 402 -1941 410
rect -1933 402 -1925 410
rect -1920 402 -1912 410
rect -1904 402 -1896 410
rect -1872 402 -1864 410
rect -1856 402 -1848 410
rect -1606 402 -1598 410
rect -1591 402 -1583 410
rect -1568 402 -1560 410
rect -857 623 -849 631
rect -842 623 -834 631
rect -825 623 -817 631
rect -809 623 -801 631
rect -794 623 -786 631
rect -781 623 -773 631
rect -766 623 -758 631
rect -748 623 -740 631
rect -733 623 -725 631
rect -716 623 -708 631
rect -701 623 -693 631
rect -688 623 -680 631
rect -673 623 -665 631
rect -649 623 -641 631
rect -633 623 -625 631
rect -618 623 -610 631
rect -605 623 -597 631
rect -590 623 -582 631
rect -571 623 -563 631
rect -555 623 -547 631
rect -525 623 -517 631
rect -508 623 -500 631
rect -495 623 -487 631
rect -480 623 -472 631
rect -374 623 -366 631
rect -359 623 -351 631
rect -342 623 -334 631
rect -327 623 -319 631
rect -314 623 -306 631
rect -299 623 -291 631
rect -275 623 -267 631
rect -259 623 -251 631
rect -244 623 -236 631
rect -231 623 -223 631
rect -216 623 -208 631
rect -174 623 -166 631
rect -158 623 -150 631
rect -143 623 -135 631
rect -126 623 -118 631
rect -113 623 -105 631
rect -98 623 -90 631
rect -60 623 -52 631
rect -44 623 -36 631
rect -29 623 -21 631
rect -16 623 -8 631
rect -1 623 7 631
rect 19 623 27 631
rect 34 623 42 631
rect 51 623 59 631
rect 64 623 72 631
rect 79 623 87 631
rect -1552 402 -1544 410
rect -1539 402 -1531 410
rect -1523 402 -1515 410
rect -1491 402 -1483 410
rect -1475 402 -1467 410
rect -1170 402 -1162 410
rect -1155 402 -1147 410
rect -1132 402 -1124 410
rect -1116 402 -1108 410
rect -1103 402 -1095 410
rect -1087 402 -1079 410
rect -1055 402 -1047 410
rect -1039 402 -1031 410
rect -662 402 -654 410
rect -647 402 -639 410
rect -624 402 -616 410
rect -608 402 -600 410
rect -595 402 -587 410
rect -579 402 -571 410
rect -547 402 -539 410
rect -531 402 -523 410
rect -318 402 -310 410
rect -303 402 -295 410
rect -280 402 -272 410
rect -264 402 -256 410
rect -251 402 -243 410
rect -235 402 -227 410
rect -203 402 -195 410
rect -187 402 -179 410
rect -60 402 -52 410
rect -45 402 -37 410
rect -22 402 -14 410
rect -6 402 2 410
rect 7 402 15 410
rect 23 402 31 410
rect 55 402 63 410
rect 71 402 79 410
<< polysilicon >>
rect -2765 949 -2762 953
rect -2723 949 -2720 953
rect -2694 949 -2691 953
rect -2678 949 -2675 953
rect -2662 949 -2659 953
rect -2645 949 -2642 953
rect -2609 949 -2606 953
rect -2593 949 -2590 953
rect -2565 949 -2562 953
rect -2312 949 -2309 953
rect -2270 949 -2267 953
rect -2241 949 -2238 953
rect -2225 949 -2222 953
rect -2209 949 -2206 953
rect -2192 949 -2189 953
rect -2156 949 -2153 953
rect -2140 949 -2137 953
rect -2112 949 -2109 953
rect -2021 949 -2018 953
rect -1979 949 -1976 953
rect -1950 949 -1947 953
rect -1934 949 -1931 953
rect -1918 949 -1915 953
rect -1901 949 -1898 953
rect -1865 949 -1862 953
rect -1849 949 -1846 953
rect -1821 949 -1818 953
rect -1778 949 -1775 953
rect -1736 949 -1733 953
rect -1707 949 -1704 953
rect -1691 949 -1688 953
rect -1675 949 -1672 953
rect -1658 949 -1655 953
rect -1622 949 -1619 953
rect -1606 949 -1603 953
rect -1578 949 -1575 953
rect -1096 949 -1093 953
rect -1054 949 -1051 953
rect -1025 949 -1022 953
rect -1009 949 -1006 953
rect -993 949 -990 953
rect -976 949 -973 953
rect -940 949 -937 953
rect -924 949 -921 953
rect -896 949 -893 953
rect -643 949 -640 953
rect -601 949 -598 953
rect -572 949 -569 953
rect -556 949 -553 953
rect -540 949 -537 953
rect -523 949 -520 953
rect -487 949 -484 953
rect -471 949 -468 953
rect -443 949 -440 953
rect -352 949 -349 953
rect -310 949 -307 953
rect -281 949 -278 953
rect -265 949 -262 953
rect -249 949 -246 953
rect -232 949 -229 953
rect -196 949 -193 953
rect -180 949 -177 953
rect -152 949 -149 953
rect -109 949 -106 953
rect -67 949 -64 953
rect -38 949 -35 953
rect -22 949 -19 953
rect -6 949 -3 953
rect 11 949 14 953
rect 47 949 50 953
rect 63 949 66 953
rect 91 949 94 953
rect -2765 819 -2762 933
rect -2723 839 -2720 933
rect -2694 839 -2691 933
rect -2723 836 -2691 839
rect -2723 818 -2720 836
rect -2694 830 -2691 836
rect -2678 830 -2675 933
rect -2662 830 -2659 933
rect -2645 830 -2642 933
rect -2765 800 -2762 811
rect -2694 817 -2691 822
rect -2678 817 -2675 822
rect -2662 817 -2659 822
rect -2723 806 -2720 810
rect -2645 800 -2642 822
rect -2765 797 -2642 800
rect -3087 617 -3084 771
rect -3070 617 -3067 741
rect -3054 617 -3051 713
rect -3038 617 -3035 688
rect -3022 617 -3019 645
rect -2994 617 -2991 621
rect -2959 617 -2956 755
rect -2943 617 -2940 741
rect -2927 617 -2924 713
rect -2911 617 -2908 688
rect -2883 617 -2880 621
rect -2850 617 -2847 727
rect -2834 617 -2831 713
rect -2818 617 -2815 688
rect -2790 617 -2787 621
rect -2751 617 -2748 700
rect -2735 617 -2732 688
rect -2624 680 -2621 857
rect -2609 804 -2606 933
rect -2593 804 -2590 933
rect -2565 804 -2562 933
rect -2609 792 -2606 796
rect -2593 792 -2590 796
rect -2565 792 -2562 796
rect -2707 617 -2704 621
rect -2673 617 -2670 622
rect -2657 617 -2654 622
rect -2641 617 -2638 622
rect -2625 617 -2622 622
rect -2610 617 -2607 675
rect -2553 667 -2552 675
rect -2544 666 -2541 909
rect -2312 819 -2309 933
rect -2270 839 -2267 933
rect -2241 839 -2238 933
rect -2270 836 -2238 839
rect -2270 818 -2267 836
rect -2241 830 -2238 836
rect -2225 830 -2222 933
rect -2209 830 -2206 933
rect -2192 830 -2189 933
rect -2312 800 -2309 811
rect -2241 817 -2238 822
rect -2225 817 -2222 822
rect -2209 817 -2206 822
rect -2270 806 -2267 810
rect -2192 800 -2189 822
rect -2312 797 -2189 800
rect -2582 617 -2579 621
rect -2516 617 -2513 770
rect -2500 617 -2497 741
rect -2484 617 -2481 713
rect -2468 617 -2465 645
rect -2440 617 -2437 621
rect -2407 617 -2404 713
rect -2391 617 -2388 755
rect -2375 617 -2372 742
rect -2347 617 -2344 621
rect -2308 617 -2305 727
rect -2292 617 -2289 713
rect -2171 705 -2168 860
rect -2156 804 -2153 933
rect -2140 804 -2137 933
rect -2112 804 -2109 933
rect -2156 792 -2153 796
rect -2140 792 -2137 796
rect -2112 792 -2109 796
rect -2091 652 -2088 909
rect -2021 819 -2018 933
rect -1979 839 -1976 933
rect -1950 839 -1947 933
rect -1979 836 -1947 839
rect -1979 818 -1976 836
rect -1950 830 -1947 836
rect -1934 830 -1931 933
rect -1918 830 -1915 933
rect -1901 830 -1898 933
rect -2021 800 -2018 811
rect -1950 817 -1947 822
rect -1934 817 -1931 822
rect -1918 817 -1915 822
rect -1979 806 -1976 810
rect -1901 800 -1898 822
rect -2021 797 -1898 800
rect -2182 649 -2088 652
rect -2264 617 -2261 621
rect -2230 617 -2227 622
rect -2214 617 -2211 622
rect -2198 617 -2195 622
rect -2182 617 -2179 649
rect -2154 617 -2151 621
rect -2033 617 -2030 741
rect -2017 617 -2014 770
rect -2001 617 -1998 645
rect -1973 617 -1970 621
rect -1934 617 -1931 755
rect -1918 617 -1915 741
rect -1880 733 -1877 862
rect -1865 804 -1862 933
rect -1849 804 -1846 933
rect -1821 804 -1818 933
rect -1865 792 -1862 796
rect -1849 792 -1846 796
rect -1821 792 -1818 796
rect -1890 617 -1887 621
rect -1833 617 -1830 622
rect -1817 617 -1814 622
rect -1800 617 -1797 911
rect -1778 819 -1775 933
rect -1736 839 -1733 933
rect -1707 839 -1704 933
rect -1736 836 -1704 839
rect -1736 818 -1733 836
rect -1707 830 -1704 836
rect -1691 830 -1688 933
rect -1675 830 -1672 933
rect -1658 830 -1655 933
rect -1778 800 -1775 811
rect -1707 817 -1704 822
rect -1691 817 -1688 822
rect -1675 817 -1672 822
rect -1736 806 -1733 810
rect -1658 800 -1655 822
rect -1778 797 -1655 800
rect -1772 617 -1769 621
rect -1653 615 -1650 645
rect -1637 615 -1634 875
rect -1622 804 -1619 933
rect -1606 804 -1603 933
rect -1578 804 -1575 933
rect -1622 792 -1619 796
rect -1606 792 -1603 796
rect -1578 792 -1575 796
rect -1609 615 -1606 619
rect -1574 615 -1571 620
rect -1557 615 -1554 909
rect -1096 819 -1093 933
rect -1054 839 -1051 933
rect -1025 839 -1022 933
rect -1054 836 -1022 839
rect -1054 818 -1051 836
rect -1025 830 -1022 836
rect -1009 830 -1006 933
rect -993 830 -990 933
rect -976 830 -973 933
rect -1096 800 -1093 811
rect -1025 817 -1022 822
rect -1009 817 -1006 822
rect -993 817 -990 822
rect -1054 806 -1051 810
rect -976 800 -973 822
rect -1096 797 -973 800
rect -1529 615 -1526 619
rect -1483 615 -1480 768
rect -1466 615 -1463 739
rect -1450 615 -1447 711
rect -1434 615 -1431 686
rect -1418 615 -1415 643
rect -1390 615 -1387 619
rect -1355 615 -1352 753
rect -1339 615 -1336 739
rect -1323 615 -1320 711
rect -1307 615 -1304 686
rect -1279 615 -1276 619
rect -1246 615 -1243 725
rect -1230 615 -1227 711
rect -1214 615 -1211 686
rect -1186 615 -1183 619
rect -1147 615 -1144 698
rect -1131 615 -1128 686
rect -955 678 -952 875
rect -940 804 -937 933
rect -924 804 -921 933
rect -896 804 -893 933
rect -940 792 -937 796
rect -924 792 -921 796
rect -896 792 -893 796
rect -1103 615 -1100 619
rect -1069 615 -1066 620
rect -1053 615 -1050 620
rect -1037 615 -1034 620
rect -1021 615 -1018 620
rect -1006 615 -1003 673
rect -875 664 -872 909
rect -643 819 -640 933
rect -601 839 -598 933
rect -572 839 -569 933
rect -601 836 -569 839
rect -601 818 -598 836
rect -572 830 -569 836
rect -556 830 -553 933
rect -540 830 -537 933
rect -523 830 -520 933
rect -643 800 -640 811
rect -572 817 -569 822
rect -556 817 -553 822
rect -540 817 -537 822
rect -601 806 -598 810
rect -523 800 -520 822
rect -643 797 -520 800
rect -978 615 -975 619
rect -3087 491 -3084 601
rect -3070 491 -3067 601
rect -3054 491 -3051 601
rect -3038 491 -3035 601
rect -3022 491 -3019 601
rect -2994 491 -2991 601
rect -2959 491 -2956 601
rect -2943 491 -2940 601
rect -2927 491 -2924 601
rect -2911 491 -2908 601
rect -2883 491 -2880 601
rect -2850 491 -2847 601
rect -2834 491 -2831 601
rect -2818 491 -2815 601
rect -2790 491 -2787 601
rect -2751 491 -2748 601
rect -2735 491 -2732 601
rect -2707 491 -2704 601
rect -2673 491 -2670 601
rect -2657 491 -2654 601
rect -2641 491 -2638 601
rect -2625 491 -2622 601
rect -2610 491 -2607 601
rect -2582 491 -2579 601
rect -2516 491 -2513 601
rect -2500 491 -2497 601
rect -2484 491 -2481 601
rect -2468 491 -2465 601
rect -2440 491 -2437 601
rect -2407 491 -2404 601
rect -2391 491 -2388 601
rect -2375 491 -2372 601
rect -2347 491 -2344 601
rect -2308 491 -2305 601
rect -2292 491 -2289 601
rect -2264 491 -2261 601
rect -2230 491 -2227 601
rect -2214 491 -2211 601
rect -2198 491 -2195 601
rect -2182 491 -2179 601
rect -2154 491 -2151 601
rect -3087 479 -3084 483
rect -3070 479 -3067 483
rect -3054 479 -3051 483
rect -3038 479 -3035 483
rect -3022 479 -3019 483
rect -2994 479 -2991 483
rect -2959 470 -2956 483
rect -2943 470 -2940 483
rect -2927 470 -2924 483
rect -2911 415 -2908 483
rect -2883 470 -2880 483
rect -2850 479 -2847 483
rect -2834 470 -2831 483
rect -2818 470 -2815 483
rect -2790 479 -2787 483
rect -2751 470 -2748 483
rect -2735 479 -2732 483
rect -2707 470 -2704 483
rect -2673 479 -2670 483
rect -2657 479 -2654 483
rect -2641 479 -2638 483
rect -2625 479 -2622 483
rect -2610 470 -2607 483
rect -2582 479 -2579 483
rect -2516 468 -2513 483
rect -2500 469 -2497 483
rect -2484 470 -2481 483
rect -2468 479 -2465 483
rect -2440 479 -2437 483
rect -2911 412 -2826 415
rect -2829 394 -2826 412
rect -2790 394 -2787 433
rect -2407 415 -2404 483
rect -2391 469 -2388 483
rect -2375 479 -2372 483
rect -2347 479 -2344 483
rect -2308 469 -2305 483
rect -2292 479 -2289 483
rect -2264 470 -2261 483
rect -2230 479 -2227 483
rect -2214 479 -2211 483
rect -2198 479 -2195 483
rect -2182 469 -2179 483
rect -2154 479 -2151 483
rect -2407 412 -2318 415
rect -2761 393 -2758 397
rect -2745 393 -2742 397
rect -2729 393 -2726 397
rect -2713 393 -2710 397
rect -2321 394 -2318 412
rect -2282 394 -2279 452
rect -2129 422 -2126 578
rect -2033 491 -2030 601
rect -2017 491 -2014 601
rect -2001 491 -1998 601
rect -1973 491 -1970 601
rect -1934 491 -1931 601
rect -1918 491 -1915 601
rect -1890 491 -1887 601
rect -1833 491 -1830 601
rect -1817 491 -1814 601
rect -1800 491 -1797 601
rect -1772 491 -1769 601
rect -2033 415 -2030 483
rect -2017 469 -2014 483
rect -2001 479 -1998 483
rect -1973 479 -1970 483
rect -1934 469 -1931 483
rect -1918 479 -1915 483
rect -1890 470 -1887 483
rect -1833 479 -1830 483
rect -1817 479 -1814 483
rect -1800 469 -1797 483
rect -1772 479 -1769 483
rect -1744 439 -1741 579
rect -1653 489 -1650 599
rect -1637 489 -1634 599
rect -1609 489 -1606 599
rect -1574 489 -1571 599
rect -1557 489 -1554 599
rect -1529 489 -1526 599
rect -2033 412 -1974 415
rect -2829 282 -2826 378
rect -2790 302 -2787 378
rect -2253 393 -2250 397
rect -2237 393 -2234 397
rect -2221 393 -2218 397
rect -2205 393 -2202 397
rect -1977 394 -1974 412
rect -1938 394 -1935 432
rect -1653 415 -1650 481
rect -1637 443 -1634 481
rect -1609 477 -1606 481
rect -1574 477 -1571 481
rect -1557 467 -1554 481
rect -1529 477 -1526 481
rect -1637 439 -1554 443
rect -1653 412 -1593 415
rect -2761 302 -2758 377
rect -2790 299 -2758 302
rect -2790 281 -2787 299
rect -2761 293 -2758 299
rect -2745 293 -2742 377
rect -2729 293 -2726 377
rect -2713 293 -2710 377
rect -2829 263 -2826 274
rect -2761 280 -2758 285
rect -2745 280 -2742 285
rect -2729 280 -2726 285
rect -2790 269 -2787 273
rect -2713 263 -2710 285
rect -2321 282 -2318 378
rect -2282 302 -2279 378
rect -1909 393 -1906 397
rect -1893 393 -1890 397
rect -1877 393 -1874 397
rect -1861 393 -1858 397
rect -1596 394 -1593 412
rect -1557 394 -1554 439
rect -1508 419 -1505 580
rect -1483 489 -1480 599
rect -1466 489 -1463 599
rect -1450 489 -1447 599
rect -1434 489 -1431 599
rect -1418 489 -1415 599
rect -1390 489 -1387 599
rect -1355 489 -1352 599
rect -1339 489 -1336 599
rect -1323 489 -1320 599
rect -1307 489 -1304 599
rect -1279 489 -1276 599
rect -1246 489 -1243 599
rect -1230 489 -1227 599
rect -1214 489 -1211 599
rect -1186 489 -1183 599
rect -1147 489 -1144 599
rect -1131 489 -1128 599
rect -1103 489 -1100 599
rect -1069 489 -1066 599
rect -1053 489 -1050 599
rect -1037 489 -1034 599
rect -1021 489 -1018 599
rect -1006 489 -1003 599
rect -978 489 -975 599
rect -953 568 -950 660
rect -847 615 -844 768
rect -831 615 -828 739
rect -815 615 -812 711
rect -799 615 -796 643
rect -771 615 -768 619
rect -738 615 -735 753
rect -722 615 -719 739
rect -706 615 -703 711
rect -678 615 -675 619
rect -639 615 -636 725
rect -623 615 -620 711
rect -502 703 -499 875
rect -487 804 -484 933
rect -471 804 -468 933
rect -443 804 -440 933
rect -487 792 -484 796
rect -471 792 -468 796
rect -443 792 -440 796
rect -422 650 -419 909
rect -352 819 -349 933
rect -310 839 -307 933
rect -281 839 -278 933
rect -310 836 -278 839
rect -310 818 -307 836
rect -281 830 -278 836
rect -265 830 -262 933
rect -249 830 -246 933
rect -232 830 -229 933
rect -352 800 -349 811
rect -281 817 -278 822
rect -265 817 -262 822
rect -249 817 -246 822
rect -310 806 -307 810
rect -232 800 -229 822
rect -352 797 -229 800
rect -513 647 -419 650
rect -595 615 -592 619
rect -561 615 -558 620
rect -545 615 -542 620
rect -529 615 -526 620
rect -513 615 -510 647
rect -485 615 -482 619
rect -364 615 -361 739
rect -348 615 -345 768
rect -332 615 -329 643
rect -304 615 -301 619
rect -265 615 -262 753
rect -249 615 -246 739
rect -211 731 -208 875
rect -196 804 -193 933
rect -180 804 -177 933
rect -152 804 -149 933
rect -196 792 -193 796
rect -180 792 -177 796
rect -152 792 -149 796
rect -221 615 -218 619
rect -164 615 -161 620
rect -148 615 -145 620
rect -131 615 -128 911
rect -109 819 -106 933
rect -67 839 -64 933
rect -38 839 -35 933
rect -67 836 -35 839
rect -67 818 -64 836
rect -38 830 -35 836
rect -22 830 -19 933
rect -6 830 -3 933
rect 11 830 14 933
rect -109 800 -106 811
rect -38 817 -35 822
rect -22 817 -19 822
rect -6 817 -3 822
rect -67 806 -64 810
rect 11 800 14 822
rect -109 797 14 800
rect 32 733 35 866
rect 47 804 50 933
rect 63 804 66 933
rect 91 804 94 933
rect 47 792 50 796
rect 63 792 66 796
rect 91 792 94 796
rect 112 740 115 909
rect -34 730 35 733
rect 46 736 115 740
rect -103 615 -100 619
rect -50 615 -47 643
rect -34 615 -31 730
rect -6 615 -3 619
rect 29 615 32 620
rect 46 615 49 736
rect 74 615 77 619
rect -847 489 -844 599
rect -831 489 -828 599
rect -815 489 -812 599
rect -799 489 -796 599
rect -771 489 -768 599
rect -738 489 -735 599
rect -722 489 -719 599
rect -706 489 -703 599
rect -678 489 -675 599
rect -639 489 -636 599
rect -623 489 -620 599
rect -595 489 -592 599
rect -561 489 -558 599
rect -545 489 -542 599
rect -529 489 -526 599
rect -513 489 -510 599
rect -485 489 -482 599
rect -1483 466 -1480 481
rect -1466 466 -1463 481
rect -1450 467 -1447 481
rect -1434 468 -1431 481
rect -1418 477 -1415 481
rect -1390 477 -1387 481
rect -1355 466 -1352 481
rect -1339 467 -1336 481
rect -1323 468 -1320 481
rect -1307 477 -1304 481
rect -1279 477 -1276 481
rect -1246 467 -1243 481
rect -1230 467 -1227 481
rect -1214 415 -1211 481
rect -1186 477 -1183 481
rect -1147 467 -1144 481
rect -1131 477 -1128 481
rect -1103 468 -1100 481
rect -1069 477 -1066 481
rect -1053 477 -1050 481
rect -1037 477 -1034 481
rect -1021 477 -1018 481
rect -1006 467 -1003 481
rect -978 477 -975 481
rect -847 466 -844 481
rect -831 467 -828 481
rect -815 468 -812 481
rect -799 477 -796 481
rect -771 477 -768 481
rect -738 477 -735 481
rect -722 467 -719 481
rect -1214 412 -1157 415
rect -2253 302 -2250 377
rect -2282 299 -2250 302
rect -2282 281 -2279 299
rect -2253 293 -2250 299
rect -2237 293 -2234 377
rect -2221 293 -2218 377
rect -2205 293 -2202 377
rect -2829 260 -2710 263
rect -2321 263 -2318 274
rect -2253 280 -2250 285
rect -2237 280 -2234 285
rect -2221 280 -2218 285
rect -2282 269 -2279 273
rect -2205 263 -2202 285
rect -1977 282 -1974 378
rect -1938 302 -1935 378
rect -1528 393 -1525 397
rect -1512 393 -1509 397
rect -1496 393 -1493 397
rect -1480 393 -1477 397
rect -1160 394 -1157 412
rect -1121 394 -1118 433
rect -706 415 -703 481
rect -678 477 -675 481
rect -639 467 -636 481
rect -623 477 -620 481
rect -595 468 -592 481
rect -561 477 -558 481
rect -545 477 -542 481
rect -529 477 -526 481
rect -513 467 -510 481
rect -485 477 -482 481
rect -706 412 -649 415
rect -1909 302 -1906 377
rect -1938 299 -1906 302
rect -1938 281 -1935 299
rect -1909 293 -1906 299
rect -1893 293 -1890 377
rect -1877 293 -1874 377
rect -1861 293 -1858 377
rect -2321 260 -2202 263
rect -1977 263 -1974 274
rect -1909 280 -1906 285
rect -1893 280 -1890 285
rect -1877 280 -1874 285
rect -1938 269 -1935 273
rect -1861 263 -1858 285
rect -1596 282 -1593 378
rect -1557 302 -1554 378
rect -1092 393 -1089 397
rect -1076 393 -1073 397
rect -1060 393 -1057 397
rect -1044 393 -1041 397
rect -652 394 -649 412
rect -613 394 -610 450
rect -460 422 -457 579
rect -364 489 -361 599
rect -348 489 -345 599
rect -332 489 -329 599
rect -304 489 -301 599
rect -265 489 -262 599
rect -249 489 -246 599
rect -221 489 -218 599
rect -164 489 -161 599
rect -148 489 -145 599
rect -131 489 -128 599
rect -103 489 -100 599
rect -364 415 -361 481
rect -348 467 -345 481
rect -332 477 -329 481
rect -304 477 -301 481
rect -265 467 -262 481
rect -249 477 -246 481
rect -221 468 -218 481
rect -164 477 -161 481
rect -148 477 -145 481
rect -131 467 -128 481
rect -103 477 -100 481
rect -75 437 -72 577
rect -50 489 -47 599
rect -34 489 -31 599
rect -6 489 -3 599
rect 29 489 32 599
rect 46 489 49 599
rect 74 489 77 599
rect -364 412 -305 415
rect -1528 302 -1525 377
rect -1557 299 -1525 302
rect -1557 281 -1554 299
rect -1528 293 -1525 299
rect -1512 293 -1509 377
rect -1496 293 -1493 377
rect -1480 293 -1477 377
rect -1977 260 -1858 263
rect -1596 263 -1593 274
rect -1528 280 -1525 285
rect -1512 280 -1509 285
rect -1496 280 -1493 285
rect -1557 269 -1554 273
rect -1480 263 -1477 285
rect -1160 282 -1157 378
rect -1121 302 -1118 378
rect -584 393 -581 397
rect -568 393 -565 397
rect -552 393 -549 397
rect -536 393 -533 397
rect -308 394 -305 412
rect -269 394 -266 432
rect -1092 302 -1089 377
rect -1121 299 -1089 302
rect -1121 281 -1118 299
rect -1092 293 -1089 299
rect -1076 293 -1073 377
rect -1060 293 -1057 377
rect -1044 293 -1041 377
rect -1596 260 -1477 263
rect -1160 263 -1157 274
rect -1092 280 -1089 285
rect -1076 280 -1073 285
rect -1060 280 -1057 285
rect -1121 269 -1118 273
rect -1044 263 -1041 285
rect -652 282 -649 378
rect -613 302 -610 378
rect -240 393 -237 397
rect -224 393 -221 397
rect -208 393 -205 397
rect -192 393 -189 397
rect -50 394 -47 481
rect -34 439 -31 481
rect -6 477 -3 481
rect 29 477 32 481
rect 46 477 49 481
rect 74 477 77 481
rect 95 449 98 580
rect 84 446 98 449
rect -34 436 -8 439
rect -11 394 -8 436
rect 84 421 87 446
rect -584 302 -581 377
rect -613 299 -581 302
rect -613 281 -610 299
rect -584 293 -581 299
rect -568 293 -565 377
rect -552 293 -549 377
rect -536 293 -533 377
rect -1160 260 -1041 263
rect -652 263 -649 274
rect -584 280 -581 285
rect -568 280 -565 285
rect -552 280 -549 285
rect -613 269 -610 273
rect -536 263 -533 285
rect -308 282 -305 378
rect -269 302 -266 378
rect 18 393 21 397
rect 34 393 37 397
rect 50 393 53 397
rect 66 393 69 397
rect -240 302 -237 377
rect -269 299 -237 302
rect -269 281 -266 299
rect -240 293 -237 299
rect -224 293 -221 377
rect -208 293 -205 377
rect -192 293 -189 377
rect -652 260 -533 263
rect -308 263 -305 274
rect -240 280 -237 285
rect -224 280 -221 285
rect -208 280 -205 285
rect -269 269 -266 273
rect -192 263 -189 285
rect -50 282 -47 378
rect -11 302 -8 378
rect 18 302 21 377
rect -11 299 21 302
rect -11 281 -8 299
rect 18 293 21 299
rect 34 293 37 377
rect 50 293 53 377
rect 66 293 69 377
rect -308 260 -189 263
rect -50 263 -47 274
rect 18 280 21 285
rect 34 280 37 285
rect 50 280 53 285
rect -11 269 -8 273
rect 66 263 69 285
rect -50 260 69 263
<< polycontact >>
rect -2773 891 -2765 899
rect -2731 878 -2723 886
rect -2686 861 -2678 869
rect -2670 848 -2662 856
rect -2617 891 -2609 899
rect -2632 849 -2624 857
rect -3084 762 -3076 770
rect -3067 733 -3059 741
rect -3051 705 -3043 713
rect -3035 680 -3027 688
rect -3019 637 -3011 645
rect -2956 747 -2947 755
rect -2940 733 -2931 741
rect -2924 705 -2916 713
rect -2908 680 -2900 688
rect -2847 719 -2839 727
rect -2831 705 -2823 713
rect -2759 692 -2751 700
rect -2815 680 -2807 688
rect -2732 680 -2724 688
rect -2632 680 -2624 688
rect -2601 878 -2593 886
rect -2573 917 -2565 925
rect -2552 901 -2544 909
rect -2607 667 -2599 675
rect -2552 667 -2544 675
rect -2320 891 -2312 899
rect -2278 878 -2270 886
rect -2233 861 -2225 869
rect -2217 848 -2209 856
rect -2164 891 -2156 899
rect -2179 851 -2171 859
rect -2513 762 -2505 770
rect -2497 733 -2489 741
rect -2481 705 -2473 713
rect -2465 637 -2457 645
rect -2404 705 -2396 713
rect -2388 747 -2380 755
rect -2372 733 -2364 741
rect -2305 719 -2297 727
rect -2289 705 -2280 713
rect -2179 705 -2171 713
rect -2148 878 -2140 886
rect -2120 917 -2112 925
rect -2099 901 -2091 909
rect -2099 692 -2091 700
rect -2029 891 -2021 899
rect -1987 878 -1979 886
rect -1942 861 -1934 869
rect -1926 848 -1918 856
rect -1873 891 -1865 899
rect -1888 851 -1880 859
rect -2030 733 -2022 741
rect -2014 762 -2006 770
rect -1998 637 -1990 645
rect -1931 747 -1923 755
rect -1915 733 -1907 741
rect -1888 733 -1880 741
rect -1857 878 -1849 886
rect -1829 917 -1821 925
rect -1808 903 -1800 911
rect -1808 719 -1800 727
rect -1786 891 -1778 899
rect -1744 878 -1736 886
rect -1699 861 -1691 869
rect -1683 848 -1675 856
rect -1630 891 -1622 899
rect -1645 848 -1637 856
rect -1645 762 -1637 770
rect -1650 637 -1642 645
rect -1614 878 -1606 886
rect -1586 917 -1578 925
rect -1565 901 -1557 909
rect -1565 747 -1557 755
rect -1104 891 -1096 899
rect -1062 878 -1054 886
rect -1017 861 -1009 869
rect -1001 848 -993 856
rect -948 891 -940 899
rect -963 852 -955 860
rect -1480 760 -1472 768
rect -1463 731 -1455 739
rect -1447 703 -1439 711
rect -1431 678 -1423 686
rect -1415 635 -1407 643
rect -1352 745 -1344 753
rect -1336 731 -1327 739
rect -1320 703 -1311 711
rect -1304 678 -1295 686
rect -1243 717 -1234 725
rect -1227 703 -1218 711
rect -1156 690 -1147 698
rect -1211 678 -1202 686
rect -1128 678 -1119 686
rect -963 678 -955 686
rect -932 878 -924 886
rect -904 917 -896 925
rect -883 901 -875 909
rect -1003 665 -995 673
rect -884 665 -875 673
rect -651 891 -643 899
rect -609 878 -601 886
rect -564 861 -556 869
rect -548 848 -540 856
rect -495 891 -487 899
rect -510 856 -502 864
rect -961 652 -953 660
rect -3002 585 -2994 593
rect -2891 585 -2883 593
rect -2798 585 -2790 593
rect -2715 585 -2707 593
rect -2681 585 -2673 593
rect -2665 573 -2657 581
rect -2649 554 -2641 562
rect -2633 537 -2625 545
rect -2590 495 -2582 503
rect -2448 585 -2440 593
rect -2355 585 -2347 593
rect -2272 585 -2264 593
rect -2238 585 -2230 593
rect -2222 573 -2214 581
rect -2206 554 -2198 562
rect -2162 495 -2154 503
rect -2137 570 -2129 578
rect -2787 422 -2779 430
rect -2279 441 -2271 449
rect -2137 422 -2129 430
rect -1981 585 -1973 593
rect -1898 585 -1890 593
rect -1841 585 -1833 593
rect -1825 573 -1817 581
rect -1780 495 -1772 503
rect -1752 571 -1744 579
rect -1752 441 -1744 449
rect -1617 583 -1609 591
rect -1582 583 -1574 591
rect -1537 572 -1529 580
rect -1516 572 -1508 580
rect -1935 421 -1927 429
rect -2753 339 -2745 347
rect -2737 311 -2729 319
rect -1516 421 -1508 429
rect -1398 583 -1390 591
rect -1287 583 -1279 591
rect -1194 583 -1186 591
rect -1111 583 -1103 591
rect -1077 583 -1069 591
rect -1061 571 -1053 579
rect -1045 552 -1037 560
rect -1029 535 -1021 543
rect -986 493 -978 501
rect -961 568 -953 576
rect -844 760 -836 768
rect -828 731 -820 739
rect -812 703 -804 711
rect -796 635 -788 643
rect -735 745 -727 753
rect -719 731 -711 739
rect -703 703 -695 711
rect -636 717 -628 725
rect -620 703 -611 711
rect -510 703 -502 711
rect -479 878 -471 886
rect -451 917 -443 925
rect -430 901 -422 909
rect -430 690 -422 698
rect -360 891 -352 899
rect -318 878 -310 886
rect -273 861 -265 869
rect -257 848 -249 856
rect -204 891 -196 899
rect -219 852 -211 860
rect -361 731 -353 739
rect -345 760 -337 768
rect -329 635 -321 643
rect -262 745 -254 753
rect -246 731 -238 739
rect -219 731 -211 739
rect -188 878 -180 886
rect -160 917 -152 925
rect -139 903 -131 911
rect -139 717 -131 725
rect -117 891 -109 899
rect -75 878 -67 886
rect -30 861 -22 869
rect -14 848 -6 856
rect 39 891 47 899
rect 24 852 32 860
rect 24 760 32 768
rect 55 878 63 886
rect 83 917 91 925
rect 104 901 112 909
rect 104 745 112 753
rect -47 635 -39 643
rect -779 583 -771 591
rect -686 583 -678 591
rect -603 583 -595 591
rect -569 583 -561 591
rect -553 571 -545 579
rect -537 552 -529 560
rect -493 493 -485 501
rect -468 568 -460 576
rect -2245 339 -2237 347
rect -2229 311 -2221 319
rect -1118 422 -1110 430
rect -1901 339 -1893 347
rect -1885 311 -1877 319
rect -610 439 -602 447
rect -468 422 -460 430
rect -312 583 -304 591
rect -229 583 -221 591
rect -172 583 -164 591
rect -156 571 -148 579
rect -111 493 -103 501
rect -83 569 -75 577
rect -83 439 -75 447
rect -14 583 -6 591
rect 21 583 29 591
rect 66 572 74 580
rect 87 572 95 580
rect -1520 339 -1512 347
rect -1504 311 -1496 319
rect -266 421 -258 429
rect -1084 339 -1076 347
rect -1068 311 -1060 319
rect 76 421 84 429
rect -576 339 -568 347
rect -560 311 -552 319
rect -232 339 -224 347
rect -216 311 -208 319
rect 26 339 34 347
rect 42 311 50 319
<< metal1 >>
rect -2783 957 -2774 965
rect -2766 957 -2761 965
rect -2753 957 -2734 965
rect -2726 957 -2718 965
rect -2710 957 -2705 965
rect -2697 957 -2689 965
rect -2681 957 -2656 965
rect -2648 957 -2640 965
rect -2632 957 -2618 965
rect -2610 957 -2603 965
rect -2595 957 -2588 965
rect -2580 957 -2575 965
rect -2567 957 -2560 965
rect -2552 957 -2321 965
rect -2313 957 -2308 965
rect -2300 957 -2281 965
rect -2273 957 -2265 965
rect -2257 957 -2252 965
rect -2244 957 -2236 965
rect -2228 957 -2203 965
rect -2195 957 -2187 965
rect -2179 957 -2165 965
rect -2157 957 -2150 965
rect -2142 957 -2135 965
rect -2127 957 -2122 965
rect -2114 957 -2107 965
rect -2099 957 -2030 965
rect -2022 957 -2017 965
rect -2009 957 -1990 965
rect -1982 957 -1974 965
rect -1966 957 -1961 965
rect -1953 957 -1945 965
rect -1937 957 -1912 965
rect -1904 957 -1896 965
rect -1888 957 -1874 965
rect -1866 957 -1859 965
rect -1851 957 -1844 965
rect -1836 957 -1831 965
rect -1823 957 -1816 965
rect -1808 957 -1787 965
rect -1779 957 -1774 965
rect -1766 957 -1747 965
rect -1739 957 -1731 965
rect -1723 957 -1718 965
rect -1710 957 -1702 965
rect -1694 957 -1669 965
rect -1661 957 -1653 965
rect -1645 957 -1631 965
rect -1623 957 -1616 965
rect -1608 957 -1601 965
rect -1593 957 -1588 965
rect -1580 957 -1573 965
rect -1565 957 -1105 965
rect -1097 957 -1092 965
rect -1084 957 -1065 965
rect -1057 957 -1049 965
rect -1041 957 -1036 965
rect -1028 957 -1020 965
rect -1012 957 -987 965
rect -979 957 -971 965
rect -963 957 -949 965
rect -941 957 -934 965
rect -926 957 -919 965
rect -911 957 -906 965
rect -898 957 -891 965
rect -883 958 -652 965
rect -883 957 -670 958
rect -654 957 -652 958
rect -644 957 -639 965
rect -631 957 -612 965
rect -604 957 -596 965
rect -588 957 -583 965
rect -575 957 -567 965
rect -559 957 -534 965
rect -526 957 -518 965
rect -510 957 -496 965
rect -488 957 -481 965
rect -473 957 -466 965
rect -458 957 -453 965
rect -445 957 -438 965
rect -430 957 -361 965
rect -353 957 -348 965
rect -340 957 -321 965
rect -313 957 -305 965
rect -297 957 -292 965
rect -284 957 -276 965
rect -268 957 -243 965
rect -235 957 -227 965
rect -219 957 -205 965
rect -197 957 -190 965
rect -182 957 -175 965
rect -167 957 -162 965
rect -154 957 -147 965
rect -139 957 -118 965
rect -110 957 -105 965
rect -97 957 -78 965
rect -70 957 -62 965
rect -54 957 -49 965
rect -41 957 -33 965
rect -25 957 0 965
rect 8 957 16 965
rect 24 957 38 965
rect 46 957 53 965
rect 61 957 68 965
rect 76 957 81 965
rect 89 957 96 965
rect 104 957 124 965
rect -2774 949 -2766 957
rect -2734 949 -2726 957
rect -2673 949 -2665 957
rect -2618 949 -2610 957
rect -2588 949 -2580 957
rect -2776 891 -2773 899
rect -2761 819 -2753 933
rect -2734 878 -2731 886
rect -2718 869 -2710 933
rect -2705 915 -2697 933
rect -2689 928 -2681 933
rect -2656 928 -2648 933
rect -2689 920 -2648 928
rect -2575 949 -2567 957
rect -2321 949 -2313 957
rect -2281 949 -2273 957
rect -2220 949 -2212 957
rect -2165 949 -2157 957
rect -2135 949 -2127 957
rect -2640 915 -2632 933
rect -2603 925 -2595 933
rect -2603 917 -2573 925
rect -2705 906 -2632 915
rect -2718 861 -2686 869
rect -2718 818 -2710 861
rect -2680 856 -2662 857
rect -2680 848 -2670 856
rect -2640 843 -2632 906
rect -2620 891 -2617 899
rect -2618 878 -2601 886
rect -2689 834 -2632 843
rect -2689 830 -2681 834
rect -2774 791 -2766 811
rect -2704 813 -2696 822
rect -2734 791 -2726 810
rect -2655 791 -2647 822
rect -2640 814 -2632 822
rect -2640 804 -2632 805
rect -2588 804 -2580 917
rect -2560 804 -2552 933
rect -2323 891 -2320 899
rect -2308 819 -2300 933
rect -2281 878 -2278 886
rect -2265 869 -2257 933
rect -2252 915 -2244 933
rect -2236 928 -2228 933
rect -2203 928 -2195 933
rect -2236 920 -2195 928
rect -2122 949 -2114 957
rect -2030 949 -2022 957
rect -1990 949 -1982 957
rect -1929 949 -1921 957
rect -1874 949 -1866 957
rect -1844 949 -1836 957
rect -2187 915 -2179 933
rect -2150 925 -2142 933
rect -2150 917 -2120 925
rect -2252 906 -2179 915
rect -2265 861 -2233 869
rect -2265 818 -2257 861
rect -2227 856 -2209 857
rect -2227 848 -2217 856
rect -2187 843 -2179 906
rect -2167 891 -2164 899
rect -2165 878 -2148 886
rect -2236 834 -2179 843
rect -2236 830 -2228 834
rect -2619 791 -2611 796
rect -2575 791 -2567 796
rect -2321 791 -2313 811
rect -2251 813 -2243 822
rect -2281 791 -2273 810
rect -2202 791 -2194 822
rect -2187 814 -2179 822
rect -2187 804 -2179 805
rect -2135 804 -2127 917
rect -2107 804 -2099 933
rect -2032 891 -2029 899
rect -2017 819 -2009 933
rect -1990 878 -1987 886
rect -1974 869 -1966 933
rect -1961 915 -1953 933
rect -1945 928 -1937 933
rect -1912 928 -1904 933
rect -1945 920 -1904 928
rect -1831 949 -1823 957
rect -1787 949 -1779 957
rect -1747 949 -1739 957
rect -1686 949 -1678 957
rect -1631 949 -1623 957
rect -1601 949 -1593 957
rect -1896 915 -1888 933
rect -1859 925 -1851 933
rect -1859 917 -1829 925
rect -1961 906 -1888 915
rect -1974 861 -1942 869
rect -1974 818 -1966 861
rect -1936 856 -1918 857
rect -1936 848 -1926 856
rect -1896 843 -1888 906
rect -1876 891 -1873 899
rect -1874 878 -1857 886
rect -1945 834 -1888 843
rect -1945 830 -1937 834
rect -2166 791 -2158 796
rect -2122 791 -2114 796
rect -2030 791 -2022 811
rect -1960 813 -1952 822
rect -1990 791 -1982 810
rect -1911 791 -1903 822
rect -1896 814 -1888 822
rect -1896 804 -1888 805
rect -1844 804 -1836 917
rect -1816 804 -1808 933
rect -1789 891 -1786 899
rect -1774 819 -1766 933
rect -1747 878 -1744 886
rect -1731 869 -1723 933
rect -1718 915 -1710 933
rect -1702 928 -1694 933
rect -1669 928 -1661 933
rect -1702 920 -1661 928
rect -1588 949 -1580 957
rect -1105 949 -1097 957
rect -1065 949 -1057 957
rect -1004 949 -996 957
rect -949 949 -941 957
rect -919 949 -911 957
rect -1653 915 -1645 933
rect -1616 925 -1608 933
rect -1616 917 -1586 925
rect -1718 906 -1645 915
rect -1731 861 -1699 869
rect -1731 818 -1723 861
rect -1693 856 -1675 857
rect -1693 848 -1683 856
rect -1653 843 -1645 906
rect -1633 891 -1630 899
rect -1631 878 -1614 886
rect -1702 834 -1645 843
rect -1702 830 -1694 834
rect -1875 791 -1867 796
rect -1831 791 -1823 796
rect -1787 791 -1779 811
rect -1717 813 -1709 822
rect -1747 791 -1739 810
rect -1668 791 -1660 822
rect -1653 814 -1645 822
rect -1653 804 -1645 805
rect -1601 804 -1593 917
rect -1573 804 -1565 933
rect -1107 891 -1104 899
rect -1092 819 -1084 933
rect -1065 878 -1062 886
rect -1049 869 -1041 933
rect -1036 915 -1028 933
rect -1020 928 -1012 933
rect -987 928 -979 933
rect -1020 920 -979 928
rect -906 949 -898 957
rect -652 949 -644 957
rect -612 949 -604 957
rect -551 949 -543 957
rect -496 949 -488 957
rect -466 949 -458 957
rect -971 915 -963 933
rect -934 925 -926 933
rect -934 917 -904 925
rect -1036 906 -963 915
rect -1049 861 -1017 869
rect -1049 818 -1041 861
rect -1011 856 -993 857
rect -1011 848 -1001 856
rect -971 843 -963 906
rect -951 891 -948 899
rect -949 878 -932 886
rect -1020 834 -963 843
rect -1020 830 -1012 834
rect -1632 791 -1624 796
rect -1588 791 -1580 796
rect -1105 791 -1097 811
rect -1035 813 -1027 822
rect -1065 791 -1057 810
rect -986 791 -978 822
rect -971 814 -963 822
rect -971 804 -963 805
rect -919 804 -911 917
rect -891 804 -883 933
rect -654 891 -651 899
rect -639 819 -631 933
rect -612 878 -609 886
rect -596 869 -588 933
rect -583 915 -575 933
rect -567 928 -559 933
rect -534 928 -526 933
rect -567 920 -526 928
rect -453 949 -445 957
rect -361 949 -353 957
rect -321 949 -313 957
rect -260 949 -252 957
rect -205 949 -197 957
rect -175 949 -167 957
rect -518 915 -510 933
rect -481 925 -473 933
rect -481 917 -451 925
rect -583 906 -510 915
rect -596 861 -564 869
rect -596 818 -588 861
rect -558 856 -540 857
rect -558 848 -548 856
rect -518 843 -510 906
rect -498 891 -495 899
rect -496 878 -479 886
rect -567 834 -510 843
rect -567 830 -559 834
rect -950 791 -942 796
rect -906 791 -898 796
rect -652 791 -644 811
rect -582 813 -574 822
rect -612 791 -604 810
rect -533 791 -525 822
rect -518 814 -510 822
rect -518 804 -510 805
rect -466 804 -458 917
rect -438 804 -430 933
rect -363 891 -360 899
rect -348 819 -340 933
rect -321 878 -318 886
rect -305 869 -297 933
rect -292 915 -284 933
rect -276 928 -268 933
rect -243 928 -235 933
rect -276 920 -235 928
rect -162 949 -154 957
rect -118 949 -110 957
rect -78 949 -70 957
rect -17 949 -9 957
rect 38 949 46 957
rect 68 949 76 957
rect -227 915 -219 933
rect -190 925 -182 933
rect -190 917 -160 925
rect -292 906 -219 915
rect -305 861 -273 869
rect -305 818 -297 861
rect -267 856 -249 857
rect -267 848 -257 856
rect -227 843 -219 906
rect -207 891 -204 899
rect -205 878 -188 886
rect -276 834 -219 843
rect -276 830 -268 834
rect -497 791 -489 796
rect -453 791 -445 796
rect -361 791 -353 811
rect -291 813 -283 822
rect -321 791 -313 810
rect -242 791 -234 822
rect -227 814 -219 822
rect -227 804 -219 805
rect -175 804 -167 917
rect -147 804 -139 933
rect -120 891 -117 899
rect -105 819 -97 933
rect -78 878 -75 886
rect -62 869 -54 933
rect -49 915 -41 933
rect -33 928 -25 933
rect 0 928 8 933
rect -33 920 8 928
rect 81 949 89 957
rect 16 915 24 933
rect 53 925 61 933
rect 53 917 83 925
rect -49 906 24 915
rect -62 861 -30 869
rect -62 818 -54 861
rect -24 856 -6 857
rect -24 848 -14 856
rect 16 843 24 906
rect 36 891 39 899
rect 38 878 55 886
rect -33 834 24 843
rect -33 830 -25 834
rect -206 791 -198 796
rect -162 791 -154 796
rect -118 791 -110 811
rect -48 813 -40 822
rect -78 791 -70 810
rect 1 791 9 822
rect 16 814 24 822
rect 16 804 24 805
rect 68 804 76 917
rect 96 804 104 933
rect 37 791 45 796
rect 81 791 89 796
rect -3116 783 -2774 791
rect -2766 783 -2760 791
rect -2752 783 -2734 791
rect -2726 783 -2717 791
rect -2709 783 -2704 791
rect -2696 783 -2687 791
rect -2679 783 -2655 791
rect -2647 783 -2638 791
rect -2630 783 -2619 791
rect -2611 783 -2603 791
rect -2595 783 -2588 791
rect -2580 783 -2575 791
rect -2567 783 -2560 791
rect -2552 783 -2321 791
rect -2313 783 -2307 791
rect -2299 783 -2281 791
rect -2273 783 -2264 791
rect -2256 783 -2251 791
rect -2243 783 -2234 791
rect -2226 783 -2202 791
rect -2194 783 -2185 791
rect -2177 783 -2166 791
rect -2158 783 -2150 791
rect -2142 783 -2135 791
rect -2127 783 -2122 791
rect -2114 783 -2107 791
rect -2099 783 -2030 791
rect -2022 783 -2016 791
rect -2008 783 -1990 791
rect -1982 783 -1973 791
rect -1965 783 -1960 791
rect -1952 783 -1943 791
rect -1935 783 -1911 791
rect -1903 783 -1894 791
rect -1886 783 -1875 791
rect -1867 783 -1859 791
rect -1851 783 -1844 791
rect -1836 783 -1831 791
rect -1823 783 -1816 791
rect -1808 783 -1787 791
rect -1779 783 -1773 791
rect -1765 783 -1747 791
rect -1739 783 -1730 791
rect -1722 783 -1717 791
rect -1709 783 -1700 791
rect -1692 783 -1668 791
rect -1660 783 -1651 791
rect -1643 783 -1632 791
rect -1624 783 -1616 791
rect -1608 783 -1601 791
rect -1593 783 -1588 791
rect -1580 783 -1573 791
rect -1565 783 -1105 791
rect -1097 783 -1091 791
rect -1083 783 -1065 791
rect -1057 783 -1048 791
rect -1040 783 -1035 791
rect -1027 783 -1018 791
rect -1010 783 -986 791
rect -978 783 -969 791
rect -961 783 -950 791
rect -942 783 -934 791
rect -926 783 -919 791
rect -911 783 -906 791
rect -898 783 -891 791
rect -883 783 -652 791
rect -644 783 -638 791
rect -630 783 -612 791
rect -604 783 -595 791
rect -587 783 -582 791
rect -574 783 -565 791
rect -557 783 -533 791
rect -525 783 -516 791
rect -508 783 -497 791
rect -489 783 -481 791
rect -473 783 -466 791
rect -458 783 -453 791
rect -445 783 -438 791
rect -430 783 -361 791
rect -353 783 -347 791
rect -339 783 -321 791
rect -313 783 -304 791
rect -296 783 -291 791
rect -283 783 -274 791
rect -266 783 -242 791
rect -234 783 -225 791
rect -217 783 -206 791
rect -198 783 -190 791
rect -182 783 -175 791
rect -167 783 -162 791
rect -154 783 -147 791
rect -139 783 -118 791
rect -110 783 -104 791
rect -96 783 -78 791
rect -70 783 -61 791
rect -53 783 -48 791
rect -40 783 -31 791
rect -23 783 1 791
rect 9 783 18 791
rect 26 783 37 791
rect 45 783 53 791
rect 61 783 68 791
rect 76 783 81 791
rect 89 783 96 791
rect 104 783 110 791
rect -3116 478 -3108 783
rect -3087 762 -3084 770
rect -3076 762 -2513 770
rect -2505 762 -2014 770
rect -2006 762 -1645 770
rect -1483 760 -1480 768
rect -1472 760 -844 768
rect -836 760 -345 768
rect -337 760 24 768
rect -3087 747 -2956 755
rect -2947 747 -2388 755
rect -2380 747 -1931 755
rect -1923 747 -1565 755
rect -1344 745 -735 753
rect -727 745 -262 753
rect -254 745 104 753
rect -3087 733 -3067 741
rect -3059 733 -2940 741
rect -2931 733 -2497 741
rect -2489 733 -2372 741
rect -2364 733 -2030 741
rect -2022 733 -1915 741
rect -1907 733 -1888 741
rect -1483 731 -1463 739
rect -1455 731 -1336 739
rect -1327 731 -828 739
rect -820 731 -719 739
rect -711 731 -361 739
rect -353 731 -246 739
rect -238 731 -219 739
rect -3087 719 -2847 727
rect -2839 719 -2305 727
rect -2297 719 -1808 727
rect -1483 717 -1243 725
rect -1234 717 -636 725
rect -628 717 -139 725
rect -3087 705 -3051 713
rect -3043 705 -2924 713
rect -2916 705 -2831 713
rect -2823 705 -2481 713
rect -2473 705 -2404 713
rect -2396 705 -2289 713
rect -2280 705 -2179 713
rect -1483 703 -1447 711
rect -1439 703 -1320 711
rect -1311 703 -1227 711
rect -1218 703 -812 711
rect -804 703 -703 711
rect -695 703 -620 711
rect -611 703 -510 711
rect -3087 692 -2759 700
rect -2751 692 -2099 700
rect -1483 690 -1156 698
rect -1147 690 -430 698
rect -3027 680 -2908 688
rect -2900 680 -2815 688
rect -2807 680 -2732 688
rect -2724 680 -2632 688
rect -1483 678 -1431 686
rect -1423 678 -1304 686
rect -1295 678 -1211 686
rect -1202 678 -1128 686
rect -1119 678 -963 686
rect -2599 667 -2552 675
rect -995 665 -884 673
rect -1520 652 -961 660
rect -1520 645 -1513 652
rect -3011 637 -2465 645
rect -2457 637 -1998 645
rect -1990 637 -1650 645
rect -1642 637 -1513 645
rect -1407 635 -796 643
rect -788 635 -329 643
rect -321 635 -47 643
rect -39 635 -20 643
rect -3103 625 -3097 633
rect -3089 625 -3080 633
rect -3072 625 -3065 633
rect -3057 625 -3048 633
rect -3040 625 -3032 633
rect -3024 625 -3017 633
rect -3009 625 -3004 633
rect -2996 625 -2989 633
rect -2981 625 -2969 633
rect -2961 625 -2954 633
rect -2946 625 -2937 633
rect -2929 625 -2921 633
rect -2913 625 -2906 633
rect -2898 625 -2893 633
rect -2885 625 -2878 633
rect -2870 625 -2860 633
rect -2852 625 -2845 633
rect -2837 625 -2828 633
rect -2820 625 -2813 633
rect -2805 625 -2800 633
rect -2792 625 -2785 633
rect -2777 625 -2761 633
rect -2753 625 -2745 633
rect -2737 625 -2730 633
rect -2722 625 -2717 633
rect -2709 625 -2702 633
rect -2694 625 -2683 633
rect -2675 625 -2667 633
rect -2659 625 -2636 633
rect -2628 625 -2621 633
rect -2613 625 -2605 633
rect -2597 625 -2592 633
rect -2584 625 -2577 633
rect -2569 625 -2526 633
rect -2518 625 -2511 633
rect -2503 625 -2494 633
rect -2486 625 -2478 633
rect -2470 625 -2463 633
rect -2455 625 -2450 633
rect -2442 625 -2435 633
rect -2427 625 -2417 633
rect -2409 625 -2402 633
rect -2394 625 -2385 633
rect -2377 625 -2370 633
rect -2362 625 -2357 633
rect -2349 625 -2342 633
rect -2334 625 -2318 633
rect -2310 625 -2302 633
rect -2294 625 -2287 633
rect -2279 625 -2274 633
rect -2266 625 -2259 633
rect -2251 625 -2240 633
rect -2232 625 -2224 633
rect -2216 625 -2194 633
rect -2186 625 -2177 633
rect -2169 625 -2164 633
rect -2156 625 -2149 633
rect -2141 625 -2043 633
rect -2035 625 -2028 633
rect -2020 625 -2011 633
rect -2003 625 -1996 633
rect -1988 625 -1983 633
rect -1975 625 -1968 633
rect -1960 625 -1944 633
rect -1936 625 -1928 633
rect -1920 625 -1913 633
rect -1905 625 -1900 633
rect -1892 625 -1885 633
rect -1877 625 -1843 633
rect -1835 625 -1827 633
rect -1819 625 -1812 633
rect -1804 625 -1795 633
rect -1787 625 -1782 633
rect -1774 625 -1767 633
rect -1759 631 -1667 633
rect 117 631 124 957
rect -1759 625 -1663 631
rect -3097 617 -3089 625
rect -3065 617 -3057 625
rect -3032 617 -3024 625
rect -3004 617 -2996 625
rect -2954 617 -2946 625
rect -2921 617 -2913 625
rect -2893 617 -2885 625
rect -2845 617 -2837 625
rect -2813 617 -2805 625
rect -3080 593 -3072 601
rect -3048 593 -3040 601
rect -3017 593 -3009 601
rect -3097 585 -3002 593
rect -3017 491 -3009 585
rect -2989 545 -2981 601
rect -2969 593 -2961 601
rect -2937 593 -2929 601
rect -2906 593 -2898 601
rect -2969 585 -2891 593
rect -2989 537 -2978 545
rect -2989 491 -2981 537
rect -2906 491 -2898 585
rect -2878 562 -2870 601
rect -2800 617 -2792 625
rect -2761 617 -2753 625
rect -2730 617 -2722 625
rect -2717 617 -2709 625
rect -2683 617 -2675 625
rect -2592 617 -2584 625
rect -2511 617 -2503 625
rect -2478 617 -2470 625
rect -2450 617 -2442 625
rect -2402 617 -2394 625
rect -2370 617 -2362 625
rect -2860 593 -2852 601
rect -2828 593 -2820 601
rect -2860 585 -2798 593
rect -2878 554 -2866 562
rect -2878 491 -2870 554
rect -2813 491 -2805 585
rect -2785 581 -2777 601
rect -2745 593 -2737 601
rect -2702 593 -2694 601
rect -2745 585 -2715 593
rect -2702 585 -2681 593
rect -2785 573 -2771 581
rect -2785 491 -2777 573
rect -2730 491 -2722 585
rect -2702 491 -2694 585
rect -2681 573 -2665 581
rect -2681 554 -2649 562
rect -2681 537 -2633 545
rect -2605 503 -2597 601
rect -2577 578 -2569 601
rect -2526 593 -2518 601
rect -2494 593 -2486 601
rect -2463 593 -2455 601
rect -2526 585 -2448 593
rect -2577 570 -2567 578
rect -2683 495 -2590 503
rect -2683 491 -2675 495
rect -2651 491 -2643 495
rect -2620 491 -2612 495
rect -2577 491 -2569 570
rect -2463 491 -2455 585
rect -2435 562 -2427 601
rect -2357 617 -2349 625
rect -2318 617 -2310 625
rect -2287 617 -2279 625
rect -2274 617 -2266 625
rect -2240 617 -2232 625
rect -2164 617 -2156 625
rect -2028 617 -2020 625
rect -1996 617 -1988 625
rect -2417 593 -2409 601
rect -2385 593 -2377 601
rect -2417 585 -2355 593
rect -2435 554 -2423 562
rect -2435 491 -2427 554
rect -2370 491 -2362 585
rect -2342 581 -2334 601
rect -2302 593 -2294 601
rect -2259 593 -2251 601
rect -2302 585 -2272 593
rect -2259 585 -2238 593
rect -2342 573 -2328 581
rect -2342 491 -2334 573
rect -2287 491 -2279 585
rect -2259 491 -2251 585
rect -2238 573 -2222 581
rect -2238 554 -2206 562
rect -2177 503 -2169 601
rect -2149 578 -2141 601
rect -1983 617 -1975 625
rect -1944 617 -1936 625
rect -1913 617 -1905 625
rect -1900 617 -1892 625
rect -1843 617 -1835 625
rect -1782 617 -1774 625
rect -1674 623 -1663 625
rect -1655 623 -1647 631
rect -1639 623 -1632 631
rect -1624 623 -1619 631
rect -1611 623 -1604 631
rect -1596 623 -1584 631
rect -1576 623 -1569 631
rect -1561 623 -1552 631
rect -1544 623 -1539 631
rect -1531 623 -1524 631
rect -1516 623 -1493 631
rect -1485 623 -1476 631
rect -1468 623 -1461 631
rect -1453 623 -1444 631
rect -1436 623 -1428 631
rect -1420 623 -1413 631
rect -1405 623 -1400 631
rect -1392 623 -1385 631
rect -1377 623 -1365 631
rect -1357 623 -1350 631
rect -1342 623 -1333 631
rect -1325 623 -1317 631
rect -1309 623 -1302 631
rect -1294 623 -1289 631
rect -1281 623 -1274 631
rect -1266 623 -1256 631
rect -1248 623 -1241 631
rect -1233 623 -1224 631
rect -1216 623 -1209 631
rect -1201 623 -1196 631
rect -1188 623 -1181 631
rect -1173 623 -1157 631
rect -1149 623 -1141 631
rect -1133 623 -1126 631
rect -1118 623 -1113 631
rect -1105 623 -1098 631
rect -1090 623 -1079 631
rect -1071 623 -1063 631
rect -1055 623 -1032 631
rect -1024 623 -1017 631
rect -1009 623 -1001 631
rect -993 623 -988 631
rect -980 623 -973 631
rect -965 623 -857 631
rect -849 623 -842 631
rect -834 623 -825 631
rect -817 623 -809 631
rect -801 623 -794 631
rect -786 623 -781 631
rect -773 623 -766 631
rect -758 623 -748 631
rect -740 623 -733 631
rect -725 623 -716 631
rect -708 623 -701 631
rect -693 623 -688 631
rect -680 623 -673 631
rect -665 623 -649 631
rect -641 623 -633 631
rect -625 623 -618 631
rect -610 623 -605 631
rect -597 623 -590 631
rect -582 623 -571 631
rect -563 623 -555 631
rect -547 623 -525 631
rect -517 623 -508 631
rect -500 623 -495 631
rect -487 623 -480 631
rect -472 623 -374 631
rect -366 623 -359 631
rect -351 623 -342 631
rect -334 623 -327 631
rect -319 623 -314 631
rect -306 623 -299 631
rect -291 623 -275 631
rect -267 623 -259 631
rect -251 623 -244 631
rect -236 623 -231 631
rect -223 623 -216 631
rect -208 623 -174 631
rect -166 623 -158 631
rect -150 623 -143 631
rect -135 623 -126 631
rect -118 623 -113 631
rect -105 623 -98 631
rect -90 623 -60 631
rect -52 623 -44 631
rect -36 623 -29 631
rect -21 623 -16 631
rect -8 623 -1 631
rect 7 623 19 631
rect 27 623 34 631
rect 42 623 51 631
rect 59 623 64 631
rect 72 623 79 631
rect 87 623 124 631
rect -2043 593 -2035 601
rect -2011 593 -2003 601
rect -2043 585 -1981 593
rect -2149 570 -2137 578
rect -3098 478 -3090 483
rect -3004 478 -2996 483
rect -2970 478 -2962 483
rect -2893 478 -2885 483
rect -2861 478 -2853 483
rect -2800 478 -2792 483
rect -2762 478 -2754 483
rect -2717 478 -2709 483
rect -2667 478 -2659 483
rect -2635 478 -2627 483
rect -2605 478 -2597 483
rect -2240 495 -2162 503
rect -2240 491 -2232 495
rect -2208 491 -2200 495
rect -2177 491 -2169 495
rect -2149 491 -2141 570
rect -1996 491 -1988 585
rect -1968 581 -1960 601
rect -1928 593 -1920 601
rect -1885 593 -1877 601
rect -1928 585 -1898 593
rect -1885 585 -1841 593
rect -1968 573 -1954 581
rect -1968 491 -1960 573
rect -1913 491 -1905 585
rect -1885 491 -1877 585
rect -1841 573 -1825 581
rect -1795 503 -1787 601
rect -1767 579 -1759 601
rect -1663 615 -1655 623
rect -1632 615 -1624 623
rect -1619 615 -1611 623
rect -1584 615 -1576 623
rect -1539 615 -1531 623
rect -1493 615 -1485 623
rect -1461 615 -1453 623
rect -1428 615 -1420 623
rect -1400 615 -1392 623
rect -1350 615 -1342 623
rect -1317 615 -1309 623
rect -1289 615 -1281 623
rect -1241 615 -1233 623
rect -1209 615 -1201 623
rect -1647 591 -1639 599
rect -1604 591 -1596 599
rect -1647 583 -1617 591
rect -1604 583 -1582 591
rect -1767 571 -1752 579
rect -1843 495 -1780 503
rect -1843 491 -1835 495
rect -1811 491 -1803 495
rect -1767 491 -1759 571
rect -2592 478 -2584 483
rect -2527 478 -2519 483
rect -2450 478 -2442 483
rect -2418 478 -2410 483
rect -2357 478 -2349 483
rect -2319 478 -2311 483
rect -2274 478 -2266 483
rect -2224 478 -2216 483
rect -2193 478 -2185 483
rect -2164 478 -2156 483
rect -2044 478 -2036 483
rect -1983 478 -1975 483
rect -1945 478 -1937 483
rect -1900 478 -1892 483
rect -1827 478 -1819 483
rect -1795 478 -1787 483
rect -1632 489 -1624 583
rect -1604 489 -1596 583
rect -1552 580 -1544 599
rect -1568 572 -1537 580
rect -1568 489 -1560 572
rect -1524 489 -1516 599
rect -1476 591 -1468 599
rect -1444 591 -1436 599
rect -1413 591 -1405 599
rect -1493 583 -1398 591
rect -1413 489 -1405 583
rect -1385 543 -1377 599
rect -1365 591 -1357 599
rect -1333 591 -1325 599
rect -1302 591 -1294 599
rect -1365 583 -1287 591
rect -1385 535 -1374 543
rect -1385 489 -1377 535
rect -1302 489 -1294 583
rect -1274 560 -1266 599
rect -1196 615 -1188 623
rect -1157 615 -1149 623
rect -1126 615 -1118 623
rect -1113 615 -1105 623
rect -1079 615 -1071 623
rect -988 615 -980 623
rect -842 615 -834 623
rect -809 615 -801 623
rect -781 615 -773 623
rect -733 615 -725 623
rect -701 615 -693 623
rect -1256 591 -1248 599
rect -1224 591 -1216 599
rect -1256 583 -1194 591
rect -1274 552 -1262 560
rect -1274 489 -1266 552
rect -1209 489 -1201 583
rect -1181 579 -1173 599
rect -1141 591 -1133 599
rect -1098 591 -1090 599
rect -1141 583 -1111 591
rect -1098 583 -1077 591
rect -1181 571 -1167 579
rect -1181 489 -1173 571
rect -1126 489 -1118 583
rect -1098 489 -1090 583
rect -1077 571 -1061 579
rect -1077 552 -1045 560
rect -1077 535 -1029 543
rect -1001 501 -993 599
rect -973 576 -965 599
rect -857 591 -849 599
rect -825 591 -817 599
rect -794 591 -786 599
rect -857 583 -779 591
rect -973 568 -961 576
rect -1782 478 -1774 483
rect -1664 478 -1656 481
rect -3116 470 -3098 478
rect -3090 470 -3081 478
rect -3073 470 -3064 478
rect -3056 470 -3048 478
rect -3040 470 -3032 478
rect -3024 470 -3017 478
rect -3009 470 -3004 478
rect -2996 470 -2989 478
rect -2981 470 -2970 478
rect -2962 470 -2953 478
rect -2945 470 -2937 478
rect -2929 470 -2921 478
rect -2913 470 -2906 478
rect -2898 470 -2893 478
rect -2885 470 -2878 478
rect -2870 470 -2861 478
rect -2853 470 -2844 478
rect -2836 470 -2828 478
rect -2820 470 -2813 478
rect -2805 470 -2800 478
rect -2792 470 -2785 478
rect -2777 470 -2762 478
rect -2754 470 -2745 478
rect -2737 470 -2730 478
rect -2722 470 -2717 478
rect -2709 470 -2702 478
rect -2694 470 -2683 478
rect -2675 470 -2667 478
rect -2659 470 -2651 478
rect -2643 470 -2635 478
rect -2627 470 -2620 478
rect -2612 470 -2605 478
rect -2597 470 -2592 478
rect -2584 470 -2577 478
rect -2569 470 -2527 478
rect -2519 470 -2510 478
rect -2502 470 -2494 478
rect -2486 470 -2478 478
rect -2470 470 -2463 478
rect -2455 470 -2450 478
rect -2442 470 -2435 478
rect -2427 470 -2418 478
rect -2410 470 -2401 478
rect -2393 470 -2385 478
rect -2377 470 -2370 478
rect -2362 470 -2357 478
rect -2349 470 -2342 478
rect -2334 470 -2319 478
rect -2311 470 -2302 478
rect -2294 470 -2287 478
rect -2279 470 -2274 478
rect -2266 470 -2259 478
rect -2251 470 -2240 478
rect -2232 470 -2224 478
rect -2216 470 -2208 478
rect -2200 470 -2193 478
rect -2185 470 -2177 478
rect -2169 470 -2164 478
rect -2156 470 -2149 478
rect -2141 470 -2044 478
rect -2036 470 -2027 478
rect -2019 470 -2011 478
rect -2003 470 -1996 478
rect -1988 470 -1983 478
rect -1975 470 -1968 478
rect -1960 470 -1945 478
rect -1937 470 -1928 478
rect -1920 470 -1913 478
rect -1905 470 -1900 478
rect -1892 470 -1885 478
rect -1877 470 -1843 478
rect -1835 470 -1827 478
rect -1819 470 -1811 478
rect -1803 470 -1795 478
rect -1787 470 -1782 478
rect -1774 470 -1767 478
rect -1759 476 -1656 478
rect -1619 476 -1611 481
rect -1584 476 -1576 481
rect -1552 476 -1544 481
rect -1079 493 -986 501
rect -1079 489 -1071 493
rect -1047 489 -1039 493
rect -1016 489 -1008 493
rect -973 489 -965 568
rect -794 489 -786 583
rect -766 560 -758 599
rect -688 615 -680 623
rect -649 615 -641 623
rect -618 615 -610 623
rect -605 615 -597 623
rect -571 615 -563 623
rect -495 615 -487 623
rect -359 615 -351 623
rect -327 615 -319 623
rect -748 591 -740 599
rect -716 591 -708 599
rect -748 583 -686 591
rect -766 552 -754 560
rect -766 489 -758 552
rect -701 489 -693 583
rect -673 579 -665 599
rect -633 591 -625 599
rect -590 591 -582 599
rect -633 583 -603 591
rect -590 583 -569 591
rect -673 571 -659 579
rect -673 489 -665 571
rect -618 489 -610 583
rect -590 489 -582 583
rect -569 571 -553 579
rect -569 552 -537 560
rect -508 501 -500 599
rect -480 576 -472 599
rect -314 615 -306 623
rect -275 615 -267 623
rect -244 615 -236 623
rect -231 615 -223 623
rect -174 615 -166 623
rect -113 615 -105 623
rect -60 615 -52 623
rect -29 615 -21 623
rect -16 615 -8 623
rect 19 615 27 623
rect 64 615 72 623
rect -374 591 -366 599
rect -342 591 -334 599
rect -374 583 -312 591
rect -480 568 -468 576
rect -1539 476 -1531 481
rect -1494 476 -1486 481
rect -1400 476 -1392 481
rect -1366 476 -1358 481
rect -1289 476 -1281 481
rect -1257 476 -1249 481
rect -1196 476 -1188 481
rect -1158 476 -1150 481
rect -1113 476 -1105 481
rect -1063 476 -1055 481
rect -1031 476 -1023 481
rect -1001 476 -993 481
rect -571 493 -493 501
rect -571 489 -563 493
rect -539 489 -531 493
rect -508 489 -500 493
rect -480 489 -472 568
rect -327 489 -319 583
rect -299 579 -291 599
rect -259 591 -251 599
rect -216 591 -208 599
rect -259 583 -229 591
rect -216 583 -172 591
rect -299 571 -285 579
rect -299 489 -291 571
rect -244 489 -236 583
rect -216 489 -208 583
rect -172 571 -156 579
rect -126 501 -118 599
rect -98 577 -90 599
rect -44 591 -36 599
rect -1 591 7 599
rect -44 583 -14 591
rect -1 583 21 591
rect -98 569 -83 577
rect -98 568 -89 569
rect -174 493 -111 501
rect -174 489 -166 493
rect -142 489 -134 493
rect -98 489 -90 568
rect -29 489 -21 583
rect -1 489 7 583
rect 51 580 59 599
rect 35 572 66 580
rect 35 489 43 572
rect 79 489 87 599
rect -988 476 -980 481
rect -858 476 -850 481
rect -781 476 -773 481
rect -749 476 -741 481
rect -688 476 -680 481
rect -650 476 -642 481
rect -605 476 -597 481
rect -555 476 -547 481
rect -524 476 -516 481
rect -495 476 -487 481
rect -375 476 -367 481
rect -314 476 -306 481
rect -276 476 -268 481
rect -231 476 -223 481
rect -158 476 -150 481
rect -126 476 -118 481
rect -113 476 -105 481
rect -61 476 -53 481
rect -16 476 -8 481
rect 19 476 27 481
rect 51 476 59 481
rect 64 476 72 481
rect -1759 470 -1664 476
rect -3116 254 -3108 470
rect -1744 468 -1664 470
rect -1656 468 -1647 476
rect -1639 468 -1632 476
rect -1624 468 -1619 476
rect -1611 468 -1604 476
rect -1596 468 -1584 476
rect -1576 468 -1568 476
rect -1560 468 -1552 476
rect -1544 468 -1539 476
rect -1531 468 -1524 476
rect -1516 468 -1494 476
rect -1486 468 -1477 476
rect -1469 468 -1460 476
rect -1452 468 -1444 476
rect -1436 468 -1428 476
rect -1420 468 -1413 476
rect -1405 468 -1400 476
rect -1392 468 -1385 476
rect -1377 468 -1366 476
rect -1358 468 -1349 476
rect -1341 468 -1333 476
rect -1325 468 -1317 476
rect -1309 468 -1302 476
rect -1294 468 -1289 476
rect -1281 468 -1274 476
rect -1266 468 -1257 476
rect -1249 468 -1240 476
rect -1232 468 -1224 476
rect -1216 468 -1209 476
rect -1201 468 -1196 476
rect -1188 468 -1181 476
rect -1173 468 -1158 476
rect -1150 468 -1141 476
rect -1133 468 -1126 476
rect -1118 468 -1113 476
rect -1105 468 -1098 476
rect -1090 468 -1079 476
rect -1071 468 -1063 476
rect -1055 468 -1047 476
rect -1039 468 -1031 476
rect -1023 468 -1016 476
rect -1008 468 -1001 476
rect -993 468 -988 476
rect -980 468 -973 476
rect -965 468 -858 476
rect -850 468 -841 476
rect -833 468 -825 476
rect -817 468 -809 476
rect -801 468 -794 476
rect -786 468 -781 476
rect -773 468 -766 476
rect -758 468 -749 476
rect -741 468 -732 476
rect -724 468 -716 476
rect -708 468 -701 476
rect -693 468 -688 476
rect -680 468 -673 476
rect -665 468 -650 476
rect -642 468 -633 476
rect -625 468 -618 476
rect -610 468 -605 476
rect -597 468 -590 476
rect -582 468 -571 476
rect -563 468 -555 476
rect -547 468 -539 476
rect -531 468 -524 476
rect -516 468 -508 476
rect -500 468 -495 476
rect -487 468 -480 476
rect -472 468 -375 476
rect -367 468 -358 476
rect -350 468 -342 476
rect -334 468 -327 476
rect -319 468 -314 476
rect -306 468 -299 476
rect -291 468 -276 476
rect -268 468 -259 476
rect -251 468 -244 476
rect -236 468 -231 476
rect -223 468 -216 476
rect -208 468 -174 476
rect -166 468 -158 476
rect -150 468 -142 476
rect -134 468 -126 476
rect -118 468 -113 476
rect -105 468 -98 476
rect -90 468 -61 476
rect -53 468 -44 476
rect -36 468 -29 476
rect -21 468 -16 476
rect -8 468 -1 476
rect 7 468 19 476
rect 27 468 35 476
rect 43 468 51 476
rect 59 468 64 476
rect 72 468 79 476
rect 87 468 88 476
rect -2271 441 -1752 449
rect -602 439 -83 447
rect -2779 422 -2137 430
rect -1927 421 -1516 429
rect -1110 422 -468 430
rect -258 421 76 429
rect 116 410 124 623
rect -2848 402 -2839 410
rect -2831 402 -2824 410
rect -2816 402 -2801 410
rect -2793 402 -2785 410
rect -2777 402 -2772 410
rect -2764 402 -2756 410
rect -2748 402 -2724 410
rect -2716 402 -2708 410
rect -2700 402 -2331 410
rect -2323 402 -2316 410
rect -2308 402 -2293 410
rect -2285 402 -2277 410
rect -2269 402 -2264 410
rect -2256 402 -2248 410
rect -2240 402 -2216 410
rect -2208 402 -2200 410
rect -2192 402 -1987 410
rect -1979 402 -1972 410
rect -1964 402 -1949 410
rect -1941 402 -1933 410
rect -1925 402 -1920 410
rect -1912 402 -1904 410
rect -1896 402 -1872 410
rect -1864 402 -1856 410
rect -1848 402 -1606 410
rect -1598 402 -1591 410
rect -1583 402 -1568 410
rect -1560 402 -1552 410
rect -1544 402 -1539 410
rect -1531 402 -1523 410
rect -1515 402 -1491 410
rect -1483 402 -1475 410
rect -1467 402 -1170 410
rect -1162 402 -1155 410
rect -1147 402 -1132 410
rect -1124 402 -1116 410
rect -1108 402 -1103 410
rect -1095 402 -1087 410
rect -1079 402 -1055 410
rect -1047 402 -1039 410
rect -1031 402 -662 410
rect -654 402 -647 410
rect -639 402 -624 410
rect -616 402 -608 410
rect -600 402 -595 410
rect -587 402 -579 410
rect -571 402 -547 410
rect -539 402 -531 410
rect -523 402 -318 410
rect -310 402 -303 410
rect -295 402 -280 410
rect -272 402 -264 410
rect -256 402 -251 410
rect -243 402 -235 410
rect -227 402 -203 410
rect -195 402 -187 410
rect -179 402 -60 410
rect -52 402 -45 410
rect -37 402 -22 410
rect -14 402 -6 410
rect 2 402 7 410
rect 15 402 23 410
rect 31 402 55 410
rect 63 402 71 410
rect 79 402 124 410
rect -2839 394 -2831 402
rect -2801 394 -2793 402
rect -2740 393 -2732 402
rect -2331 394 -2323 402
rect -2293 394 -2285 402
rect -2824 282 -2816 378
rect -2785 369 -2777 370
rect -2772 360 -2764 377
rect -2756 373 -2748 377
rect -2724 373 -2716 377
rect -2756 364 -2716 373
rect -2232 393 -2224 402
rect -1987 394 -1979 402
rect -1949 394 -1941 402
rect -2708 360 -2700 377
rect -2772 351 -2700 360
rect -2765 339 -2753 347
rect -2785 281 -2777 331
rect -2747 311 -2737 319
rect -2708 306 -2700 351
rect -2756 297 -2700 306
rect -2756 293 -2748 297
rect -2839 254 -2831 274
rect -2771 277 -2763 285
rect -2801 254 -2793 273
rect -2723 254 -2715 285
rect -2708 277 -2700 285
rect -2316 282 -2308 378
rect -2277 369 -2269 370
rect -2264 360 -2256 377
rect -2248 373 -2240 377
rect -2216 373 -2208 377
rect -2248 364 -2208 373
rect -1888 393 -1880 402
rect -1606 394 -1598 402
rect -1568 394 -1560 402
rect -2200 360 -2192 377
rect -2264 351 -2192 360
rect -2257 339 -2245 347
rect -2277 281 -2269 331
rect -2239 311 -2229 319
rect -2200 306 -2192 351
rect -2248 297 -2192 306
rect -2248 293 -2240 297
rect -2331 254 -2323 274
rect -2263 276 -2255 285
rect -2293 254 -2285 273
rect -2215 254 -2207 285
rect -2200 277 -2192 285
rect -1972 282 -1964 378
rect -1933 369 -1925 370
rect -1920 360 -1912 377
rect -1904 373 -1896 377
rect -1872 373 -1864 377
rect -1904 364 -1864 373
rect -1507 393 -1499 402
rect -1170 394 -1162 402
rect -1132 394 -1124 402
rect -1856 360 -1848 377
rect -1920 351 -1848 360
rect -1913 339 -1901 347
rect -2200 267 -2192 268
rect -1933 281 -1925 331
rect -1895 311 -1885 319
rect -1856 306 -1848 351
rect -1904 297 -1848 306
rect -1904 293 -1896 297
rect -1987 254 -1979 274
rect -1919 276 -1911 285
rect -1949 254 -1941 273
rect -1871 254 -1863 285
rect -1856 277 -1848 285
rect -1591 282 -1583 378
rect -1552 369 -1544 370
rect -1539 360 -1531 377
rect -1523 373 -1515 377
rect -1491 373 -1483 377
rect -1523 364 -1483 373
rect -1071 393 -1063 402
rect -662 394 -654 402
rect -624 394 -616 402
rect -1475 360 -1467 377
rect -1539 351 -1467 360
rect -1532 339 -1520 347
rect -1856 267 -1848 268
rect -1552 281 -1544 331
rect -1514 311 -1504 319
rect -1475 306 -1467 351
rect -1523 297 -1467 306
rect -1523 293 -1515 297
rect -1606 254 -1598 274
rect -1538 276 -1530 285
rect -1568 254 -1560 273
rect -1490 254 -1482 285
rect -1475 277 -1467 285
rect -1155 282 -1147 378
rect -1116 369 -1108 370
rect -1103 360 -1095 377
rect -1087 373 -1079 377
rect -1055 373 -1047 377
rect -1087 364 -1047 373
rect -563 393 -555 402
rect -318 394 -310 402
rect -280 394 -272 402
rect -1037 360 -1029 377
rect -1103 351 -1029 360
rect -1096 339 -1084 347
rect -1475 267 -1467 268
rect -1116 281 -1108 331
rect -1078 311 -1068 319
rect -1037 306 -1029 351
rect -1087 297 -1029 306
rect -1087 293 -1079 297
rect -1170 254 -1162 274
rect -1102 277 -1094 285
rect -1132 254 -1124 273
rect -1054 254 -1046 285
rect -1037 277 -1029 285
rect -647 282 -639 378
rect -608 369 -600 370
rect -595 360 -587 377
rect -579 373 -571 377
rect -547 373 -539 377
rect -579 364 -539 373
rect -219 393 -211 402
rect -60 394 -52 402
rect -22 394 -14 402
rect -531 360 -523 377
rect -595 351 -523 360
rect -588 339 -576 347
rect -608 281 -600 331
rect -570 311 -560 319
rect -531 306 -523 351
rect -579 297 -523 306
rect -579 293 -571 297
rect -662 254 -654 274
rect -594 277 -586 285
rect -624 254 -616 273
rect -546 254 -538 285
rect -531 277 -523 285
rect -303 282 -295 378
rect -264 369 -256 370
rect -251 360 -243 377
rect -235 373 -227 377
rect -203 373 -195 377
rect -235 364 -195 373
rect 39 393 47 402
rect -187 360 -179 377
rect -251 351 -179 360
rect -244 339 -232 347
rect -264 281 -256 331
rect -226 311 -216 319
rect -187 306 -179 351
rect -235 297 -179 306
rect -235 293 -227 297
rect -318 254 -310 274
rect -250 276 -242 285
rect -280 254 -272 273
rect -202 254 -194 285
rect -187 277 -179 285
rect -45 282 -37 378
rect -6 369 2 370
rect 7 360 15 377
rect 23 373 31 377
rect 55 373 63 377
rect 23 364 63 373
rect 71 360 79 377
rect 7 351 79 360
rect 14 339 26 347
rect -187 267 -179 268
rect -6 281 2 331
rect 32 311 42 319
rect 71 306 79 351
rect 23 297 79 306
rect 23 293 31 297
rect -60 254 -52 274
rect 8 276 16 285
rect -22 254 -14 273
rect 56 254 64 285
rect 71 277 79 285
rect 71 267 79 268
rect -3116 246 -2839 254
rect -2831 246 -2823 254
rect -2815 246 -2801 254
rect -2793 246 -2784 254
rect -2776 246 -2771 254
rect -2763 246 -2754 254
rect -2746 246 -2723 254
rect -2715 246 -2706 254
rect -2698 246 -2331 254
rect -2323 246 -2315 254
rect -2307 246 -2293 254
rect -2285 246 -2276 254
rect -2268 246 -2263 254
rect -2255 246 -2246 254
rect -2238 246 -2215 254
rect -2207 246 -2198 254
rect -2190 246 -1987 254
rect -1979 246 -1971 254
rect -1963 246 -1949 254
rect -1941 246 -1932 254
rect -1924 246 -1919 254
rect -1911 246 -1902 254
rect -1894 246 -1871 254
rect -1863 246 -1854 254
rect -1846 246 -1606 254
rect -1598 246 -1590 254
rect -1582 246 -1568 254
rect -1560 246 -1551 254
rect -1543 246 -1538 254
rect -1530 246 -1521 254
rect -1513 246 -1490 254
rect -1482 246 -1473 254
rect -1465 246 -1170 254
rect -1162 246 -1154 254
rect -1146 246 -1132 254
rect -1124 246 -1115 254
rect -1107 246 -1102 254
rect -1094 246 -1085 254
rect -1077 246 -1054 254
rect -1046 246 -1037 254
rect -1029 246 -662 254
rect -654 246 -646 254
rect -638 246 -624 254
rect -616 246 -607 254
rect -599 246 -594 254
rect -586 246 -577 254
rect -569 246 -546 254
rect -538 246 -529 254
rect -521 246 -318 254
rect -310 246 -302 254
rect -294 246 -280 254
rect -272 246 -263 254
rect -255 246 -250 254
rect -242 246 -233 254
rect -225 246 -202 254
rect -194 246 -185 254
rect -177 246 -60 254
rect -52 246 -44 254
rect -36 246 -22 254
rect -14 246 -5 254
rect 3 246 8 254
rect 16 246 25 254
rect 33 246 56 254
rect 64 246 73 254
rect 81 246 87 254
<< m2contact >>
rect -2783 891 -2776 899
rect -2742 878 -2734 886
rect -2753 848 -2745 856
rect -2689 848 -2680 857
rect -2628 891 -2620 899
rect -2626 878 -2618 886
rect -2704 804 -2696 813
rect -2640 805 -2632 814
rect -2330 891 -2323 899
rect -2289 878 -2281 886
rect -2300 848 -2292 856
rect -2236 848 -2227 857
rect -2175 891 -2167 899
rect -2173 878 -2165 886
rect -2251 804 -2243 813
rect -2187 805 -2179 814
rect -2040 891 -2032 899
rect -1998 878 -1990 886
rect -2009 848 -2001 856
rect -1945 848 -1936 857
rect -1884 891 -1876 899
rect -1882 878 -1874 886
rect -1960 804 -1952 813
rect -1896 805 -1888 814
rect -1797 891 -1789 899
rect -1755 878 -1747 886
rect -1766 848 -1758 856
rect -1702 848 -1693 857
rect -1641 891 -1633 899
rect -1639 878 -1631 886
rect -1717 804 -1709 813
rect -1653 805 -1645 814
rect -1115 891 -1107 899
rect -1073 878 -1065 886
rect -1084 848 -1076 856
rect -1020 848 -1011 857
rect -959 891 -951 899
rect -957 878 -949 886
rect -1035 804 -1027 813
rect -971 805 -963 814
rect -661 891 -654 899
rect -620 878 -612 886
rect -631 848 -623 856
rect -567 848 -558 857
rect -506 891 -498 899
rect -504 878 -496 886
rect -582 804 -574 813
rect -518 805 -510 814
rect -371 891 -363 899
rect -329 878 -321 886
rect -340 848 -332 856
rect -276 848 -267 857
rect -215 891 -207 899
rect -213 878 -205 886
rect -291 804 -283 813
rect -227 805 -219 814
rect -128 891 -120 899
rect -86 878 -78 886
rect -97 848 -89 856
rect -33 848 -24 857
rect 28 891 36 899
rect 30 878 38 886
rect -48 804 -40 813
rect 16 805 24 814
rect -2978 537 -2970 545
rect -2866 554 -2858 562
rect -2771 573 -2763 581
rect -2689 573 -2681 581
rect -2689 554 -2681 562
rect -2689 537 -2681 545
rect -2423 554 -2415 562
rect -2328 573 -2320 581
rect -2246 573 -2238 581
rect -2246 554 -2238 562
rect -1954 573 -1946 581
rect -1849 573 -1841 581
rect -1374 535 -1366 543
rect -1262 552 -1254 560
rect -1167 571 -1159 579
rect -1085 571 -1077 579
rect -1085 552 -1077 560
rect -1085 535 -1077 543
rect -754 552 -746 560
rect -659 571 -651 579
rect -577 571 -569 579
rect -577 552 -569 560
rect -285 571 -277 579
rect -180 571 -172 579
rect -2785 370 -2777 378
rect -2773 339 -2765 347
rect -2785 331 -2777 339
rect -2816 311 -2808 319
rect -2755 311 -2747 319
rect -2771 269 -2763 277
rect -2277 370 -2269 378
rect -2265 339 -2257 347
rect -2277 331 -2269 339
rect -2308 311 -2300 319
rect -2708 269 -2700 277
rect -2247 311 -2239 319
rect -2263 267 -2255 276
rect -1933 370 -1925 378
rect -1921 339 -1913 347
rect -1933 331 -1925 339
rect -1964 311 -1956 319
rect -2200 268 -2192 277
rect -1903 311 -1895 319
rect -1919 267 -1911 276
rect -1552 370 -1544 378
rect -1540 339 -1532 347
rect -1552 331 -1544 339
rect -1583 311 -1575 319
rect -1856 268 -1848 277
rect -1522 311 -1514 319
rect -1538 267 -1530 276
rect -1116 370 -1108 378
rect -1104 339 -1096 347
rect -1116 331 -1108 339
rect -1147 311 -1139 319
rect -1475 268 -1467 277
rect -1086 311 -1078 319
rect -1102 268 -1094 277
rect -608 370 -600 378
rect -596 339 -588 347
rect -608 331 -600 339
rect -639 311 -631 319
rect -1037 268 -1029 277
rect -578 311 -570 319
rect -594 268 -586 277
rect -264 370 -256 378
rect -252 339 -244 347
rect -264 331 -256 339
rect -295 311 -287 319
rect -531 268 -523 277
rect -234 311 -226 319
rect -250 267 -242 276
rect -6 370 2 378
rect 6 339 14 347
rect -6 331 2 339
rect -37 311 -29 319
rect -187 268 -179 277
rect 24 311 32 319
rect 8 267 16 276
rect 71 268 79 277
<< metal2 >>
rect -2776 891 -2628 899
rect -2323 891 -2175 899
rect -2032 891 -1884 899
rect -1789 891 -1641 899
rect -1107 891 -959 899
rect -654 891 -506 899
rect -363 891 -215 899
rect -120 891 28 899
rect -2734 878 -2626 886
rect -2281 878 -2173 886
rect -1990 878 -1882 886
rect -1747 878 -1639 886
rect -1065 878 -957 886
rect -612 878 -504 886
rect -321 878 -213 886
rect -78 878 30 886
rect -2753 856 -2689 857
rect -2745 848 -2689 856
rect -2300 856 -2236 857
rect -2292 848 -2236 856
rect -2009 856 -1945 857
rect -2001 848 -1945 856
rect -1766 856 -1702 857
rect -1758 848 -1702 856
rect -1084 856 -1020 857
rect -1076 848 -1020 856
rect -631 856 -567 857
rect -623 848 -567 856
rect -340 856 -276 857
rect -332 848 -276 856
rect -97 856 -33 857
rect -89 848 -33 856
rect -2704 813 -2640 814
rect -2696 805 -2640 813
rect -2696 804 -2632 805
rect -2251 813 -2187 814
rect -2243 805 -2187 813
rect -2243 804 -2179 805
rect -1960 813 -1896 814
rect -1952 805 -1896 813
rect -1952 804 -1888 805
rect -1717 813 -1653 814
rect -1709 805 -1653 813
rect -1709 804 -1645 805
rect -1035 813 -971 814
rect -1027 805 -971 813
rect -1027 804 -963 805
rect -582 813 -518 814
rect -574 805 -518 813
rect -574 804 -510 805
rect -291 813 -227 814
rect -283 805 -227 813
rect -283 804 -219 805
rect -48 813 16 814
rect -40 805 16 813
rect -40 804 24 805
rect -2763 573 -2689 581
rect -2320 573 -2246 581
rect -1946 573 -1849 581
rect -1159 571 -1085 579
rect -651 571 -577 579
rect -277 571 -180 579
rect -2858 554 -2689 562
rect -2415 554 -2246 562
rect -1254 552 -1085 560
rect -746 552 -577 560
rect -2970 537 -2689 545
rect -1366 535 -1085 543
rect -2785 347 -2777 370
rect -2277 347 -2269 370
rect -1933 347 -1925 370
rect -1552 347 -1544 370
rect -1116 347 -1108 370
rect -608 347 -600 370
rect -264 347 -256 370
rect -6 347 2 370
rect -2785 339 -2773 347
rect -2277 339 -2265 347
rect -1933 339 -1921 347
rect -1552 339 -1540 347
rect -1116 339 -1104 347
rect -608 339 -596 347
rect -264 339 -252 347
rect -6 339 6 347
rect -2808 311 -2755 319
rect -2300 311 -2247 319
rect -1956 311 -1903 319
rect -1575 311 -1522 319
rect -1139 311 -1086 319
rect -631 311 -578 319
rect -287 311 -234 319
rect -29 311 24 319
rect -2763 269 -2708 277
rect -2263 276 -2200 277
rect -2255 268 -2200 276
rect -2255 267 -2192 268
rect -1919 276 -1856 277
rect -1911 268 -1856 276
rect -1911 267 -1848 268
rect -1538 276 -1475 277
rect -1530 268 -1475 276
rect -1094 268 -1037 277
rect -586 268 -531 277
rect -250 276 -187 277
rect -1530 267 -1467 268
rect -242 268 -187 276
rect -242 267 -179 268
rect 8 276 71 277
rect 16 268 71 276
rect 16 267 79 268
<< labels >>
rlabel metal1 -1568 905 -1568 905 1 g4
rlabel metal1 -1649 868 -1649 868 1 p4
rlabel metal2 -1788 894 -1788 894 1 a4
rlabel metal2 -1746 881 -1746 881 1 b4
rlabel metal2 -2031 896 -2031 896 1 a5
rlabel metal2 -1989 882 -1989 882 1 b5
rlabel metal1 -1893 868 -1893 868 1 p5
rlabel metal1 -1811 907 -1811 907 1 g5
rlabel metal2 -2775 896 -2775 896 1 a7
rlabel metal2 -2733 881 -2733 881 1 b7
rlabel metal1 -2636 868 -2636 868 1 p7
rlabel metal1 -2555 907 -2555 907 1 g7
rlabel metal2 -2321 895 -2321 895 1 a6
rlabel metal2 -2280 881 -2280 881 1 b6
rlabel metal1 -2183 869 -2183 869 1 p6
rlabel metal1 -2102 906 -2102 906 1 g6
rlabel metal1 -2704 332 -2704 332 1 s7
rlabel metal1 -2196 333 -2196 333 1 s6
rlabel metal1 -1852 331 -1852 331 1 s5
rlabel metal2 -1105 894 -1105 894 1 a3
rlabel metal1 -965 868 -965 868 1 p3
rlabel metal1 -887 906 -887 906 1 g3
rlabel metal2 -1063 881 -1063 881 1 b3
rlabel metal2 -119 895 -119 895 1 a0
rlabel metal1 21 867 21 867 1 p0
rlabel metal2 -76 881 -76 881 1 b0
rlabel metal1 99 906 99 906 1 g0
rlabel metal1 -144 905 -144 905 1 g1
rlabel metal1 -224 869 -224 869 1 p1
rlabel metal2 -320 882 -320 882 1 b1
rlabel metal2 -362 894 -362 894 1 a1
rlabel metal1 -435 905 -435 905 1 g2
rlabel metal1 -514 868 -514 868 1 p2
rlabel metal2 -653 894 -653 894 1 a2
rlabel metal2 -611 882 -611 882 1 b2
rlabel metal1 -1471 332 -1471 332 1 s4
rlabel metal1 -183 328 -183 328 1 s1
rlabel metal1 -528 331 -528 331 1 s2
rlabel metal1 -94 568 -94 568 1 c2
rlabel metal1 -969 573 -969 573 1 c4
rlabel metal1 -1520 576 -1520 576 1 c5
rlabel metal1 -1762 572 -1762 572 1 c6
rlabel metal1 -2145 575 -2145 575 1 c7
rlabel metal1 -1032 330 -1032 330 1 s3
rlabel metal1 -2572 573 -2572 573 1 c8
rlabel metal1 74 328 74 328 1 s0
rlabel metal1 -21 639 -21 639 3 c0
rlabel metal1 82 563 82 563 1 c1
rlabel metal1 109 786 109 786 1 gnd
rlabel metal1 -475 568 -475 568 1 c3
rlabel metal1 108 961 108 961 5 vdd
rlabel metal1 12 587 12 587 1 and1
rlabel metal1 -203 587 -203 587 1 and2
rlabel metal1 -293 576 -293 576 1 and3
<< end >>
